module otn_frame_rom
#(
    parameter                                   NB_DATA     = 256,
    parameter                                   NB_ADDRESS  = 9
)
(
    // OUTPUTS
    output  wire    [NB_DATA-1:0]               o_data ,
    output  wire                                o_valid ,

    // INPUTS
    input   wire    [NB_ADDRESS-1:0]            i_address ,
    input   wire                                i_valid
);

    // LOCAL PARAMETERS
    localparam                                  NB_BYTE     = 8;
    localparam                                  N_ADDRESS   = 2**NB_ADDRESS;       // 2**9 = 512
    localparam                                  NB_ROW      = 4;

    // INTERNAL SIGNAL
    wire            [NB_DATA-1:0]               data    [N_ADDRESS-1:0] ;
    wire            [7*NB_BYTE-1:0]             fas ;
    wire            [7*NB_BYTE-1:0]             otu_oh ;
    wire            [2*NB_BYTE-1:0]             opu_oh ;
    wire            [14*NB_BYTE-1:0]            odu_oh ;
    wire            [8*NB_BYTE-1:0]             pl  [2*N_ADDRESS-1:0] ;
    wire            [8*NB_BYTE-1:0]             fs  [NB_ROW-1:0] ;

    assign fas      = 56'h F6F6F628282828;
    assign otu_oh   = 56'h FFFFFFFFFFFFFF;
    assign opu_oh   = 16'h AAAA;

    generate
        genvar ii;
        for( ii == 0; ii<(2*N_ADDRESS); ii=ii+1 )
        begin: begin_genfor_pl
            assign pl[ii] = { 32'd0, ii };
        end
    endgenerate

    generate
        genvar jj;
        for( jj == 0; jj<NB_ROW; jj==jj+1 )
        begin: begin_genfor_fs
            assign fs[jj] = { 8'hF5, 32'd0, jj };
        end
    endgenerate

    generate
        genvar hh;
        for( hh == 0; hh<NB_ROW-1; hh==hh+1 )
        begin: begin_genfor_fs
            assign odu_oh[hh] = { 8'h44, 72'd0, hh };
        end
    endgenerate

    assign data[0]      =   { fas,  otu_oh, opu_oh,     pl[0],      pl[1]       };      // ROW 1
    assign data[1]      =   { pl[2],        pl[3],      pl[4],      pl[5]       };
    assign data[2]      =   { pl[6],        pl[7],      pl[8],      pl[9]       };
    assign data[3]      =   { pl[10],       pl[11],     pl[12],     pl[13]      };
    assign data[4]      =   { pl[14],       pl[15],     pl[16],     pl[17]      };
    assign data[5]      =   { pl[18],       pl[19],     pl[20],     pl[21]      };
    assign data[6]      =   { pl[22],       pl[23],     pl[24],     pl[25]      };
    assign data[7]      =   { pl[26],       pl[27],     pl[28],     pl[29]      };
    assign data[8]      =   { pl[30],       pl[31],     pl[32],     pl[33]      };
    assign data[9]      =   { pl[34],       pl[35],     pl[36],     pl[37]      };
    assign data[10]     =   { pl[38],       pl[39],     pl[40],     pl[41]      };
    assign data[11]     =   { pl[42],       pl[43],     pl[44],     pl[45]      };
    assign data[12]     =   { pl[46],       pl[47],     pl[48],     pl[49]      };
    assign data[13]     =   { pl[50],       pl[51],     pl[52],     pl[53]      };
    assign data[14]     =   { pl[54],       pl[55],     pl[56],     pl[57]      };
    assign data[15]     =   { pl[58],       pl[59],     pl[60],     pl[61]      };
    assign data[16]     =   { pl[62],       pl[63],     pl[64],     pl[65]      };
    assign data[17]     =   { pl[66],       pl[67],     pl[68],     pl[69]      };
    assign data[18]     =   { pl[70],       pl[71],     pl[72],     pl[73]      };
    assign data[19]     =   { pl[74],       pl[75],     pl[76],     pl[77]      };
    assign data[20]     =   { pl[78],       pl[79],     pl[80],     pl[81]      };
    assign data[21]     =   { pl[82],       pl[83],     pl[84],     pl[85]      };
    assign data[22]     =   { pl[86],       pl[87],     pl[88],     pl[89]      };
    assign data[23]     =   { pl[90],       pl[91],     pl[92],     pl[93]      };
    assign data[24]     =   { pl[94],       pl[95],     pl[96],     pl[97]      };
    assign data[25]     =   { pl[98],       pl[99],     pl[100],    pl[101]     };
    assign data[26]     =   { pl[102],      pl[103],    pl[104],    pl[105]     };
    assign data[27]     =   { pl[106],      pl[107],    pl[108],    pl[109]     };
    assign data[28]     =   { pl[110],      pl[111],    pl[112],    pl[113]     };
    assign data[29]     =   { pl[114],      pl[115],    pl[116],    pl[117]     };
    assign data[30]     =   { pl[118],      pl[119],    pl[120],    pl[121]     };
    assign data[31]     =   { pl[122],      pl[123],    pl[124],    pl[125]     };
    assign data[32]     =   { pl[126],      pl[127],    pl[128],    pl[129]     };
    assign data[33]     =   { pl[130],      pl[131],    pl[132],    pl[133]     };
    assign data[34]     =   { pl[134],      pl[135],    pl[136],    pl[137]     };
    assign data[35]     =   { pl[138],      pl[139],    pl[140],    pl[141]     };
    assign data[36]     =   { pl[142],      pl[143],    pl[144],    pl[145]     };
    assign data[37]     =   { pl[146],      pl[147],    pl[148],    pl[149]     };
    assign data[38]     =   { pl[150],      pl[151],    pl[152],    pl[153]     };
    assign data[39]     =   { pl[154],      pl[155],    pl[156],    pl[157]     };
    assign data[40]     =   { pl[158],      pl[159],    pl[160],    pl[161]     };
    assign data[41]     =   { pl[162],      pl[163],    pl[164],    pl[165]     };
    assign data[42]     =   { pl[166],      pl[167],    pl[168],    pl[169]     };
    assign data[43]     =   { pl[170],      pl[171],    pl[172],    pl[173]     };
    assign data[44]     =   { pl[174],      pl[175],    pl[176],    pl[177]     };
    assign data[45]     =   { pl[178],      pl[179],    pl[180],    pl[181]     };
    assign data[46]     =   { pl[182],      pl[183],    pl[184],    pl[185]     };
    assign data[47]     =   { pl[186],      pl[187],    pl[188],    pl[189]     };
    assign data[48]     =   { pl[190],      pl[191],    pl[192],    pl[193]     };
    assign data[49]     =   { pl[194],      pl[195],    pl[196],    pl[197]     };
    assign data[50]     =   { pl[198],      pl[199],    pl[200],    pl[201]     };
    assign data[51]     =   { pl[202],      pl[203],    pl[204],    pl[205]     };
    assign data[52]     =   { pl[206],      pl[207],    pl[208],    pl[209]     };
    assign data[53]     =   { pl[210],      pl[211],    pl[212],    pl[213]     };
    assign data[54]     =   { pl[214],      pl[215],    pl[216],    pl[217]     };
    assign data[55]     =   { pl[218],      pl[219],    pl[220],    pl[221]     };
    assign data[56]     =   { pl[222],      pl[223],    pl[224],    pl[225]     };
    assign data[57]     =   { pl[226],      pl[227],    pl[228],    pl[229]     };
    assign data[58]     =   { pl[230],      pl[231],    pl[232],    pl[233]     };
    assign data[59]     =   { pl[234],      pl[235],    pl[236],    pl[237]     };
    assign data[60]     =   { pl[238],      pl[239],    pl[240],    pl[241]     };
    assign data[61]     =   { pl[242],      pl[243],    pl[244],    pl[245]     };
    assign data[62]     =   { pl[246],      pl[247],    pl[248],    pl[249]     };
    assign data[63]     =   { pl[250],      pl[251],    pl[252],    pl[253]     };
    assign data[64]     =   { pl[254],      pl[255],    pl[256],    pl[257]     };
    assign data[65]     =   { pl[258],      pl[259],    pl[260],    pl[261]     };
    assign data[66]     =   { pl[262],      pl[263],    pl[264],    pl[265]     };
    assign data[67]     =   { pl[266],      pl[267],    pl[268],    pl[269]     };
    assign data[68]     =   { pl[270],      pl[271],    pl[272],    pl[273]     };
    assign data[69]     =   { pl[274],      pl[275],    pl[276],    pl[277]     };
    assign data[70]     =   { pl[278],      pl[279],    pl[280],    pl[281]     };
    assign data[71]     =   { pl[282],      pl[283],    pl[284],    pl[285]     };
    assign data[72]     =   { pl[286],      pl[287],    pl[288],    pl[289]     };
    assign data[73]     =   { pl[290],      pl[291],    pl[292],    pl[293]     };
    assign data[74]     =   { pl[294],      pl[295],    pl[296],    pl[297]     };
    assign data[75]     =   { pl[298],      pl[299],    pl[300],    pl[301]     };
    assign data[76]     =   { pl[302],      pl[303],    pl[304],    pl[305]     };
    assign data[77]     =   { pl[306],      pl[307],    pl[308],    pl[309]     };
    assign data[78]     =   { pl[310],      pl[311],    pl[312],    pl[313]     };
    assign data[79]     =   { pl[314],      pl[315],    pl[316],    pl[317]     };
    assign data[80]     =   { pl[318],      pl[319],    pl[320],    pl[321]     };
    assign data[81]     =   { pl[322],      pl[323],    pl[324],    pl[325]     };
    assign data[82]     =   { pl[326],      pl[327],    pl[328],    pl[329]     };
    assign data[83]     =   { pl[330],      pl[331],    pl[332],    pl[333]     };
    assign data[84]     =   { pl[334],      pl[335],    pl[336],    pl[337]     };
    assign data[85]     =   { pl[338],      pl[339],    pl[340],    pl[341]     };
    assign data[86]     =   { pl[342],      pl[343],    pl[344],    pl[345]     };
    assign data[87]     =   { pl[346],      pl[347],    pl[348],    pl[349]     };
    assign data[88]     =   { pl[350],      pl[351],    pl[352],    pl[353]     };
    assign data[89]     =   { pl[354],      pl[355],    pl[356],    pl[357]     };
    assign data[90]     =   { pl[358],      pl[359],    pl[360],    pl[361]     };
    assign data[91]     =   { pl[362],      pl[363],    pl[364],    pl[365]     };
    assign data[92]     =   { pl[366],      pl[367],    pl[368],    pl[369]     };
    assign data[93]     =   { pl[370],      pl[371],    pl[372],    pl[373]     };
    assign data[94]     =   { pl[374],      pl[375],    pl[376],    pl[377]     };
    assign data[95]     =   { pl[378],      pl[379],    pl[380],    pl[381]     };
    assign data[96]     =   { pl[382],      pl[383],    pl[384],    pl[385]     };
    assign data[97]     =   { pl[386],      pl[387],    pl[388],    pl[389]     };
    assign data[98]     =   { pl[390],      pl[391],    pl[392],    pl[393]     };
    assign data[99]     =   { pl[394],      pl[395],    pl[396],    pl[397]     };
    assign data[100]    =   { pl[398],      pl[399],    pl[400],    pl[401]     };
    assign data[101]    =   { pl[402],      pl[403],    pl[404],    pl[405]     };
    assign data[102]    =   { pl[406],      pl[407],    pl[408],    pl[409]     };
    assign data[103]    =   { pl[410],      pl[411],    pl[412],    pl[413]     };
    assign data[104]    =   { pl[414],      pl[415],    pl[416],    pl[417]     };
    assign data[105]    =   { pl[418],      pl[419],    pl[420],    pl[421]     };
    assign data[106]    =   { pl[422],      pl[423],    pl[424],    pl[425]     };
    assign data[107]    =   { pl[426],      pl[427],    pl[428],    pl[429]     };
    assign data[108]    =   { pl[430],      pl[431],    pl[432],    pl[433]     };
    assign data[109]    =   { pl[434],      pl[435],    pl[436],    pl[437]     };
    assign data[110]    =   { pl[438],      pl[439],    pl[440],    pl[441]     };
    assign data[111]    =   { pl[442],      pl[443],    pl[444],    pl[445]     };
    assign data[112]    =   { pl[446],      pl[447],    pl[448],    pl[449]     };
    assign data[113]    =   { pl[450],      pl[451],    pl[452],    pl[453]     };
    assign data[114]    =   { pl[454],      pl[455],    pl[456],    pl[457]     };
    assign data[115]    =   { pl[458],      pl[459],    pl[460],    pl[461]     };
    assign data[116]    =   { pl[462],      pl[463],    pl[464],    pl[465]     };
    assign data[117]    =   { pl[466],      pl[467],    pl[468],    pl[469]     };
    assign data[118]    =   { pl[470],      pl[471],    pl[472],    pl[473]     };
    assign data[119]    =   { pl[474],      fs[0],      fec[0],     fec[1]      };
    assign data[120]    =   { fec[2],       fec[3],     fec[4],     fec[5]      };
    assign data[121]    =   { fec[6],       fec[7],     fec[8],     fec[9]      };
    assign data[122]    =   { fec[10],      fec[11],    fec[12],    fec[13]     };
    assign data[123]    =   { fec[14],      fec[15],    fec[16],    fec[17]     };
    assign data[124]    =   { fec[18],      fec[19],    fec[20],    fec[21]     };
    assign data[125]    =   { fec[22],      fec[23],    fec[24],    fec[25]     };
    assign data[126]    =   { fec[26],      fec[27],    fec[28],    fec[29]     };

    assign data[127]    =   { fec[30],      fec[31],    odu_oh[0],  opu_oh      };      // ROW 2
    assign data[128]    =   { pl[475],      pl[476],    pl[477],    pl[478]     };
    assign data[129]    =   { pl[479],      pl[480],    pl[481],    pl[482]     };
    assign data[130]    =   { pl[483],      pl[484],    pl[485],    pl[486]     };
    assign data[131]    =   { pl[487],      pl[488],    pl[489],    pl[490]     };
    assign data[132]    =   { pl[491],      pl[492],    pl[493],    pl[494]     };
    assign data[133]    =   { pl[495],      pl[496],    pl[497],    pl[498]     };
    assign data[134]    =   { pl[499],      pl[500],    pl[501],    pl[502]     };
    assign data[135]    =   { pl[503],      pl[504],    pl[505],    pl[506]     };
    assign data[136]    =   { pl[507],      pl[508],    pl[509],    pl[510]     };
    assign data[137]    =   { pl[511],      pl[512],    pl[513],    pl[514]     };
    assign data[138]    =   { pl[515],      pl[516],    pl[517],    pl[518]     };
    assign data[139]    =   { pl[519],      pl[520],    pl[521],    pl[522]     };
    assign data[140]    =   { pl[523],      pl[524],    pl[525],    pl[526]     };
    assign data[141]    =   { pl[527],      pl[528],    pl[529],    pl[530]     };
    assign data[142]    =   { pl[531],      pl[532],    pl[533],    pl[534]     };
    assign data[143]    =   { pl[535],      pl[536],    pl[537],    pl[538]     };
    assign data[144]    =   { pl[539],      pl[540],    pl[541],    pl[542]     };
    assign data[145]    =   { pl[543],      pl[544],    pl[545],    pl[546]     };
    assign data[146]    =   { pl[547],      pl[548],    pl[549],    pl[550]     };
    assign data[147]    =   { pl[551],      pl[552],    pl[553],    pl[554]     };
    assign data[148]    =   { pl[555],      pl[556],    pl[557],    pl[558]     };
    assign data[149]    =   { pl[559],      pl[560],    pl[561],    pl[562]     };
    assign data[150]    =   { pl[563],      pl[564],    pl[565],    pl[566]     };
    assign data[151]    =   { pl[567],      pl[568],    pl[569],    pl[570]     };
    assign data[152]    =   { pl[571],      pl[572],    pl[573],    pl[574]     };
    assign data[153]    =   { pl[575],      pl[576],    pl[577],    pl[578]     };
    assign data[154]    =   { pl[579],      pl[580],    pl[581],    pl[582]     };
    assign data[155]    =   { pl[583],      pl[584],    pl[585],    pl[586]     };
    assign data[156]    =   { pl[587],      pl[588],    pl[589],    pl[590]     };
    assign data[157]    =   { pl[591],      pl[592],    pl[593],    pl[594]     };
    assign data[158]    =   { pl[595],      pl[596],    pl[597],    pl[598]     };
    assign data[159]    =   { pl[599],      pl[600],    pl[601],    pl[602]     };
    assign data[160]    =   { pl[603],      pl[604],    pl[605],    pl[606]     };
    assign data[161]    =   { pl[607],      pl[608],    pl[609],    pl[610]     };
    assign data[162]    =   { pl[611],      pl[612],    pl[613],    pl[614]     };
    assign data[163]    =   { pl[615],      pl[616],    pl[617],    pl[618]     };
    assign data[164]    =   { pl[619],      pl[620],    pl[621],    pl[622]     };
    assign data[165]    =   { pl[623],      pl[624],    pl[625],    pl[626]     };
    assign data[166]    =   { pl[627],      pl[628],    pl[629],    pl[630]     };
    assign data[167]    =   { pl[631],      pl[632],    pl[633],    pl[634]     };
    assign data[168]    =   { pl[635],      pl[636],    pl[637],    pl[638]     };
    assign data[169]    =   { pl[639],      pl[640],    pl[641],    pl[642]     };
    assign data[170]    =   { pl[643],      pl[644],    pl[645],    pl[646]     };
    assign data[171]    =   { pl[647],      pl[648],    pl[649],    pl[650]     };
    assign data[172]    =   { pl[651],      pl[652],    pl[653],    pl[654]     };
    assign data[173]    =   { pl[655],      pl[656],    pl[657],    pl[658]     };
    assign data[174]    =   { pl[659],      pl[660],    pl[661],    pl[662]     };
    assign data[175]    =   { pl[663],      pl[664],    pl[665],    pl[666]     };
    assign data[176]    =   { pl[667],      pl[668],    pl[669],    pl[670]     };
    assign data[177]    =   { pl[671],      pl[672],    pl[673],    pl[674]     };
    assign data[178]    =   { pl[675],      pl[676],    pl[677],    pl[678]     };
    assign data[179]    =   { pl[679],      pl[680],    pl[681],    pl[682]     };
    assign data[180]    =   { pl[683],      pl[684],    pl[685],    pl[686]     };
    assign data[181]    =   { pl[687],      pl[688],    pl[689],    pl[690]     };
    assign data[182]    =   { pl[691],      pl[692],    pl[693],    pl[694]     };
    assign data[183]    =   { pl[695],      pl[696],    pl[697],    pl[698]     };
    assign data[184]    =   { pl[699],      pl[700],    pl[701],    pl[702]     };
    assign data[185]    =   { pl[703],      pl[704],    pl[705],    pl[706]     };
    assign data[186]    =   { pl[707],      pl[708],    pl[709],    pl[710]     };
    assign data[187]    =   { pl[711],      pl[712],    pl[713],    pl[714]     };
    assign data[188]    =   { pl[715],      pl[716],    pl[717],    pl[718]     };
    assign data[189]    =   { pl[719],      pl[720],    pl[721],    pl[722]     };
    assign data[190]    =   { pl[723],      pl[724],    pl[725],    pl[726]     };
    assign data[191]    =   { pl[727],      pl[728],    pl[729],    pl[730]     };
    assign data[192]    =   { pl[731],      pl[732],    pl[733],    pl[734]     };
    assign data[193]    =   { pl[735],      pl[736],    pl[737],    pl[738]     };
    assign data[194]    =   { pl[739],      pl[740],    pl[741],    pl[742]     };
    assign data[195]    =   { pl[743],      pl[744],    pl[745],    pl[746]     };
    assign data[196]    =   { pl[747],      pl[748],    pl[749],    pl[750]     };
    assign data[197]    =   { pl[751],      pl[752],    pl[753],    pl[754]     };
    assign data[198]    =   { pl[755],      pl[756],    pl[757],    pl[758]     };
    assign data[199]    =   { pl[759],      pl[760],    pl[761],    pl[762]     };
    assign data[200]    =   { pl[763],      pl[764],    pl[765],    pl[766]     };
    assign data[201]    =   { pl[767],      pl[768],    pl[769],    pl[770]     };
    assign data[202]    =   { pl[771],      pl[772],    pl[773],    pl[774]     };
    assign data[203]    =   { pl[775],      pl[776],    pl[777],    pl[778]     };
    assign data[204]    =   { pl[779],      pl[780],    pl[781],    pl[782]     };
    assign data[205]    =   { pl[783],      pl[784],    pl[785],    pl[786]     };
    assign data[206]    =   { pl[787],      pl[788],    pl[789],    pl[790]     };
    assign data[207]    =   { pl[791],      pl[792],    pl[793],    pl[794]     };
    assign data[208]    =   { pl[795],      pl[796],    pl[797],    pl[798]     };
    assign data[209]    =   { pl[799],      pl[800],    pl[801],    pl[802]     };
    assign data[210]    =   { pl[803],      pl[804],    pl[805],    pl[806]     };
    assign data[211]    =   { pl[807],      pl[808],    pl[809],    pl[810]     };
    assign data[212]    =   { pl[811],      pl[812],    pl[813],    pl[814]     };
    assign data[213]    =   { pl[815],      pl[816],    pl[817],    pl[818]     };
    assign data[214]    =   { pl[819],      pl[820],    pl[821],    pl[822]     };
    assign data[215]    =   { pl[823],      pl[824],    pl[825],    pl[826]     };
    assign data[216]    =   { pl[827],      pl[828],    pl[829],    pl[830]     };
    assign data[217]    =   { pl[831],      pl[832],    pl[833],    pl[834]     };
    assign data[218]    =   { pl[835],      pl[836],    pl[837],    pl[838]     };
    assign data[219]    =   { pl[839],      pl[840],    pl[841],    pl[842]     };
    assign data[220]    =   { pl[843],      pl[844],    pl[845],    pl[846]     };
    assign data[221]    =   { pl[847],      pl[848],    pl[849],    pl[850]     };
    assign data[222]    =   { pl[851],      pl[852],    pl[853],    pl[854]     };
    assign data[223]    =   { pl[855],      pl[856],    pl[857],    pl[858]     };
    assign data[224]    =   { pl[859],      pl[860],    pl[861],    pl[862]     };
    assign data[225]    =   { pl[863],      pl[864],    pl[865],    pl[866]     };
    assign data[226]    =   { pl[867],      pl[868],    pl[869],    pl[870]     };
    assign data[227]    =   { pl[871],      pl[872],    pl[873],    pl[874]     };
    assign data[228]    =   { pl[875],      pl[876],    pl[877],    pl[878]     };
    assign data[229]    =   { pl[879],      pl[880],    pl[881],    pl[882]     };
    assign data[230]    =   { pl[883],      pl[884],    pl[885],    pl[886]     };
    assign data[231]    =   { pl[887],      pl[888],    pl[889],    pl[890]     };
    assign data[232]    =   { pl[891],      pl[892],    pl[893],    pl[894]     };
    assign data[233]    =   { pl[895],      pl[896],    pl[897],    pl[898]     };
    assign data[234]    =   { pl[899],      pl[900],    pl[901],    pl[902]     };
    assign data[235]    =   { pl[903],      pl[904],    pl[905],    pl[906]     };
    assign data[236]    =   { pl[907],      pl[908],    pl[909],    pl[910]     };
    assign data[237]    =   { pl[911],      pl[912],    pl[913],    pl[914]     };
    assign data[238]    =   { pl[915],      pl[916],    pl[917],    pl[918]     };
    assign data[239]    =   { pl[919],      pl[920],    pl[921],    pl[922]     };
    assign data[240]    =   { pl[923],      pl[924],    pl[925],    pl[926]     };
    assign data[241]    =   { pl[927],      pl[928],    pl[929],    pl[930]     };
    assign data[242]    =   { pl[931],      pl[932],    pl[933],    pl[934]     };
    assign data[243]    =   { pl[935],      pl[936],    pl[937],    pl[938]     };
    assign data[244]    =   { pl[939],      pl[940],    pl[941],    pl[942]     };
    assign data[245]    =   { pl[943],      pl[944],    pl[945],    pl[946]     };
    assign data[246]    =   { pl[947],      pl[948],    pl[949],    fs[1]       };
    assign data[247]    =   { fec[32],      fec[33],    fec[34],    fec[35]     };
    assign data[248]    =   { fec[36],      fec[37],    fec[38],    fec[39]     };
    assign data[249]    =   { fec[40],      fec[41],    fec[42],    fec[43]     };
    assign data[250]    =   { fec[44],      fec[45],    fec[46],    fec[47]     };
    assign data[251]    =   { fec[48],      fec[49],    fec[50],    fec[51]     };
    assign data[252]    =   { fec[52],      fec[53],    fec[54],    fec[55]     };
    assign data[253]    =   { fec[56],      fec[57],    fec[58],    fec[59]     };
    assign data[254]    =   { fec[60],      fec[61],    fec[62],    fec[63]     };

    assign data[255]    =   { odu_oh[1],    opu_oh,     pl[950],    pl[951]     };      // ROW 3
    assign data[256]    =   { pl[952],      pl[953],    pl[954],    pl[955]     };
    assign data[257]    =   { pl[956],      pl[957],    pl[958],    pl[959]     };
    assign data[258]    =   { pl[960],      pl[961],    pl[962],    pl[963]     };
    assign data[259]    =   { pl[964],      pl[965],    pl[966],    pl[967]     };
    assign data[260]    =   { pl[968],      pl[969],    pl[970],    pl[971]     };
    assign data[261]    =   { pl[972],      pl[973],    pl[974],    pl[975]     };
    assign data[262]    =   { pl[976],      pl[977],    pl[978],    pl[979]     };
    assign data[263]    =   { pl[980],      pl[981],    pl[982],    pl[983]     };
    assign data[264]    =   { pl[984],      pl[985],    pl[986],    pl[987]     };
    assign data[265]    =   { pl[988],      pl[989],    pl[990],    pl[991]     };
    assign data[266]    =   { pl[992],      pl[993],    pl[994],    pl[995]     };
    assign data[267]    =   { pl[996],      pl[997],    pl[998],    pl[999]     };
    assign data[268]    =   { pl[1000],     pl[1001],   pl[1002],   pl[1003]    };
    assign data[269]    =   { pl[1004],     pl[1005],   pl[1006],   pl[1007]    };
    assign data[270]    =   { pl[1008],     pl[1009],   pl[1010],   pl[1011]    };
    assign data[271]    =   { pl[1012],     pl[1013],   pl[1014],   pl[1015]    };
    assign data[272]    =   { pl[1016],     pl[1017],   pl[1018],   pl[1019]    };
    assign data[273]    =   { pl[1020],     pl[1021],   pl[1022],   pl[1023]    };
    assign data[274]    =   { pl[1024],     pl[1025],   pl[1026],   pl[1027]    };
    assign data[275]    =   { pl[1028],     pl[1029],   pl[1030],   pl[1031]    };
    assign data[276]    =   { pl[1032],     pl[1033],   pl[1034],   pl[1035]    };
    assign data[277]    =   { pl[1036],     pl[1037],   pl[1038],   pl[1039]    };
    assign data[278]    =   { pl[1040],     pl[1041],   pl[1042],   pl[1043]    };
    assign data[279]    =   { pl[1044],     pl[1045],   pl[1046],   pl[1047]    };
    assign data[280]    =   { pl[1048],     pl[1049],   pl[1050],   pl[1051]    };
    assign data[281]    =   { pl[1052],     pl[1053],   pl[1054],   pl[1055]    };
    assign data[282]    =   { pl[1056],     pl[1057],   pl[1058],   pl[1059]    };
    assign data[283]    =   { pl[1060],     pl[1061],   pl[1062],   pl[1063]    };
    assign data[284]    =   { pl[1064],     pl[1065],   pl[1066],   pl[1067]    };
    assign data[285]    =   { pl[1068],     pl[1069],   pl[1070],   pl[1071]    };
    assign data[286]    =   { pl[1072],     pl[1073],   pl[1074],   pl[1075]    };
    assign data[287]    =   { pl[1076],     pl[1077],   pl[1078],   pl[1079]    };
    assign data[288]    =   { pl[1080],     pl[1081],   pl[1082],   pl[1083]    };
    assign data[289]    =   { pl[1084],     pl[1085],   pl[1086],   pl[1087]    };
    assign data[290]    =   { pl[1088],     pl[1089],   pl[1090],   pl[1091]    };
    assign data[291]    =   { pl[1092],     pl[1093],   pl[1094],   pl[1095]    };
    assign data[292]    =   { pl[1096],     pl[1097],   pl[1098],   pl[1099]    };
    assign data[293]    =   { pl[1100],     pl[1101],   pl[1102],   pl[1103]    };
    assign data[294]    =   { pl[1104],     pl[1105],   pl[1106],   pl[1107]    };
    assign data[295]    =   { pl[1108],     pl[1109],   pl[1110],   pl[1111]    };
    assign data[296]    =   { pl[1112],     pl[1113],   pl[1114],   pl[1115]    };
    assign data[297]    =   { pl[1116],     pl[1117],   pl[1118],   pl[1119]    };
    assign data[298]    =   { pl[1120],     pl[1121],   pl[1122],   pl[1123]    };
    assign data[299]    =   { pl[1124],     pl[1125],   pl[1126],   pl[1127]    };
    assign data[300]    =   { pl[1128],     pl[1129],   pl[1130],   pl[1131]    };
    assign data[301]    =   { pl[1132],     pl[1133],   pl[1134],   pl[1135]    };
    assign data[302]    =   { pl[1136],     pl[1137],   pl[1138],   pl[1139]    };
    assign data[303]    =   { pl[1140],     pl[1141],   pl[1142],   pl[1143]    };
    assign data[304]    =   { pl[1144],     pl[1145],   pl[1146],   pl[1147]    };
    assign data[305]    =   { pl[1148],     pl[1149],   pl[1150],   pl[1151]    };
    assign data[306]    =   { pl[1152],     pl[1153],   pl[1154],   pl[1155]    };
    assign data[307]    =   { pl[1156],     pl[1157],   pl[1158],   pl[1159]    };
    assign data[308]    =   { pl[1160],     pl[1161],   pl[1162],   pl[1163]    };
    assign data[309]    =   { pl[1164],     pl[1165],   pl[1166],   pl[1167]    };
    assign data[310]    =   { pl[1168],     pl[1169],   pl[1170],   pl[1171]    };
    assign data[311]    =   { pl[1172],     pl[1173],   pl[1174],   pl[1175]    };
    assign data[312]    =   { pl[1176],     pl[1177],   pl[1178],   pl[1179]    };
    assign data[313]    =   { pl[1180],     pl[1181],   pl[1182],   pl[1183]    };
    assign data[314]    =   { pl[1184],     pl[1185],   pl[1186],   pl[1187]    };
    assign data[315]    =   { pl[1188],     pl[1189],   pl[1190],   pl[1191]    };
    assign data[316]    =   { pl[1192],     pl[1193],   pl[1194],   pl[1195]    };
    assign data[317]    =   { pl[1196],     pl[1197],   pl[1198],   pl[1199]    };
    assign data[318]    =   { pl[1200],     pl[1201],   pl[1202],   pl[1203]    };
    assign data[319]    =   { pl[1204],     pl[1205],   pl[1206],   pl[1207]    };
    assign data[320]    =   { pl[1208],     pl[1209],   pl[1210],   pl[1211]    };
    assign data[321]    =   { pl[1212],     pl[1213],   pl[1214],   pl[1215]    };
    assign data[322]    =   { pl[1216],     pl[1217],   pl[1218],   pl[1219]    };
    assign data[323]    =   { pl[1220],     pl[1221],   pl[1222],   pl[1223]    };
    assign data[324]    =   { pl[1224],     pl[1225],   pl[1226],   pl[1227]    };
    assign data[325]    =   { pl[1228],     pl[1229],   pl[1230],   pl[1231]    };
    assign data[326]    =   { pl[1232],     pl[1233],   pl[1234],   pl[1235]    };
    assign data[327]    =   { pl[1236],     pl[1237],   pl[1238],   pl[1239]    };
    assign data[328]    =   { pl[1240],     pl[1241],   pl[1242],   pl[1243]    };
    assign data[329]    =   { pl[1244],     pl[1245],   pl[1246],   pl[1247]    };
    assign data[330]    =   { pl[1248],     pl[1249],   pl[1250],   pl[1251]    };
    assign data[331]    =   { pl[1252],     pl[1253],   pl[1254],   pl[1255]    };
    assign data[332]    =   { pl[1256],     pl[1257],   pl[1258],   pl[1259]    };
    assign data[333]    =   { pl[1260],     pl[1261],   pl[1262],   pl[1263]    };
    assign data[334]    =   { pl[1264],     pl[1265],   pl[1266],   pl[1267]    };
    assign data[335]    =   { pl[1268],     pl[1269],   pl[1270],   pl[1271]    };
    assign data[336]    =   { pl[1272],     pl[1273],   pl[1274],   pl[1275]    };
    assign data[337]    =   { pl[1276],     pl[1277],   pl[1278],   pl[1279]    };
    assign data[338]    =   { pl[1280],     pl[1281],   pl[1282],   pl[1283]    };
    assign data[339]    =   { pl[1284],     pl[1285],   pl[1286],   pl[1287]    };
    assign data[340]    =   { pl[1288],     pl[1289],   pl[1290],   pl[1291]    };
    assign data[341]    =   { pl[1292],     pl[1293],   pl[1294],   pl[1295]    };
    assign data[342]    =   { pl[1296],     pl[1297],   pl[1298],   pl[1299]    };
    assign data[343]    =   { pl[1300],     pl[1301],   pl[1302],   pl[1303]    };
    assign data[344]    =   { pl[1304],     pl[1305],   pl[1306],   pl[1307]    };
    assign data[345]    =   { pl[1308],     pl[1309],   pl[1310],   pl[1311]    };
    assign data[346]    =   { pl[1312],     pl[1313],   pl[1314],   pl[1315]    };
    assign data[347]    =   { pl[1316],     pl[1317],   pl[1318],   pl[1319]    };
    assign data[348]    =   { pl[1320],     pl[1321],   pl[1322],   pl[1323]    };
    assign data[349]    =   { pl[1324],     pl[1325],   pl[1326],   pl[1327]    };
    assign data[350]    =   { pl[1328],     pl[1329],   pl[1330],   pl[1331]    };
    assign data[351]    =   { pl[1332],     pl[1333],   pl[1334],   pl[1335]    };
    assign data[352]    =   { pl[1336],     pl[1337],   pl[1338],   pl[1339]    };
    assign data[353]    =   { pl[1340],     pl[1341],   pl[1342],   pl[1343]    };
    assign data[354]    =   { pl[1344],     pl[1345],   pl[1346],   pl[1347]    };
    assign data[355]    =   { pl[1348],     pl[1349],   pl[1350],   pl[1351]    };
    assign data[356]    =   { pl[1352],     pl[1353],   pl[1354],   pl[1355]    };
    assign data[357]    =   { pl[1356],     pl[1357],   pl[1358],   pl[1359]    };
    assign data[358]    =   { pl[1360],     pl[1361],   pl[1362],   pl[1363]    };
    assign data[359]    =   { pl[1364],     pl[1365],   pl[1366],   pl[1367]    };
    assign data[360]    =   { pl[1368],     pl[1369],   pl[1370],   pl[1371]    };
    assign data[361]    =   { pl[1372],     pl[1373],   pl[1374],   pl[1375]    };
    assign data[362]    =   { pl[1376],     pl[1377],   pl[1378],   pl[1379]    };
    assign data[363]    =   { pl[1380],     pl[1381],   pl[1382],   pl[1383]    };
    assign data[364]    =   { pl[1384],     pl[1385],   pl[1386],   pl[1387]    };
    assign data[365]    =   { pl[1388],     pl[1389],   pl[1390],   pl[1391]    };
    assign data[366]    =   { pl[1392],     pl[1393],   pl[1394],   pl[1395]    };
    assign data[367]    =   { pl[1396],     pl[1397],   pl[1398],   pl[1399]    };
    assign data[368]    =   { pl[1400],     pl[1401],   pl[1402],   pl[1403]    };
    assign data[369]    =   { pl[1404],     pl[1405],   pl[1406],   pl[1407]    };
    assign data[370]    =   { pl[1408],     pl[1409],   pl[1410],   pl[1411]    };
    assign data[371]    =   { pl[1412],     pl[1413],   pl[1414],   pl[1415]    };
    assign data[372]    =   { pl[1416],     pl[1417],   pl[1418],   pl[1419]    };
    assign data[373]    =   { pl[1420],     pl[1421],   pl[1422],   pl[1423]    };
    assign data[374]    =   { pl[1424],     fs[2],      fec[64],    fec[65]     };
    assign data[375]    =   { fec[66],      fec[67],    fec[68],    fec[69]     };
    assign data[376]    =   { fec[70],      fec[71],    fec[72],    fec[73]     };
    assign data[377]    =   { fec[74],      fec[75],    fec[76],    fec[77]     };
    assign data[378]    =   { fec[78],      fec[79],    fec[80],    fec[81]     };
    assign data[379]    =   { fec[82],      fec[83],    fec[84],    fec[85]     };
    assign data[380]    =   { fec[86],      fec[87],    fec[88],    fec[89]     };
    assign data[381]    =   { fec[90],      fec[91],    fec[92],    fec[93]     };

    assign data[382]    =   { fec[94],      fec[95],    odu_oh[2],  opu_oh      };      //ROW 4
    assign data[383]    =   { pl[1425],     pl[1426],   pl[1427],   pl[1428]    };
    assign data[384]    =   { pl[1429],     pl[1430],   pl[1431],   pl[1432]    };
    assign data[385]    =   { pl[1433],     pl[1434],   pl[1435],   pl[1436]    };
    assign data[386]    =   { pl[1437],     pl[1438],   pl[1439],   pl[1440]    };
    assign data[387]    =   { pl[1441],     pl[1442],   pl[1443],   pl[1444]    };
    assign data[388]    =   { pl[1445],     pl[1446],   pl[1447],   pl[1448]    };
    assign data[389]    =   { pl[1449],     pl[1450],   pl[1451],   pl[1452]    };
    assign data[390]    =   { pl[1453],     pl[1454],   pl[1455],   pl[1456]    };
    assign data[391]    =   { pl[1457],     pl[1458],   pl[1459],   pl[1460]    };
    assign data[392]    =   { pl[1461],     pl[1462],   pl[1463],   pl[1464]    };
    assign data[393]    =   { pl[1465],     pl[1466],   pl[1467],   pl[1468]    };
    assign data[394]    =   { pl[1469],     pl[1470],   pl[1471],   pl[1472]    };
    assign data[395]    =   { pl[1473],     pl[1474],   pl[1475],   pl[1476]    };
    assign data[396]    =   { pl[1477],     pl[1478],   pl[1479],   pl[1480]    };
    assign data[397]    =   { pl[1481],     pl[1482],   pl[1483],   pl[1484]    };
    assign data[398]    =   { pl[1485],     pl[1486],   pl[1487],   pl[1488]    };
    assign data[399]    =   { pl[1489],     pl[1490],   pl[1491],   pl[1492]    };
    assign data[400]    =   { pl[1493],     pl[1494],   pl[1495],   pl[1496]    };
    assign data[401]    =   { pl[1497],     pl[1498],   pl[1499],   pl[1500]    };
    assign data[402]    =   { pl[1501],     pl[1502],   pl[1503],   pl[1504]    };
    assign data[403]    =   { pl[1505],     pl[1506],   pl[1507],   pl[1508]    };
    assign data[404]    =   { pl[1509],     pl[1510],   pl[1511],   pl[1512]    };
    assign data[405]    =   { pl[1513],     pl[1514],   pl[1515],   pl[1516]    };
    assign data[406]    =   { pl[1517],     pl[1518],   pl[1519],   pl[1520]    };
    assign data[407]    =   { pl[1521],     pl[1522],   pl[1523],   pl[1524]    };
    assign data[408]    =   { pl[1525],     pl[1526],   pl[1527],   pl[1528]    };
    assign data[409]    =   { pl[1529],     pl[1530],   pl[1531],   pl[1532]    };
    assign data[410]    =   { pl[1533],     pl[1534],   pl[1535],   pl[1536]    };
    assign data[411]    =   { pl[1537],     pl[1538],   pl[1539],   pl[1540]    };
    assign data[412]    =   { pl[1541],     pl[1542],   pl[1543],   pl[1544]    };
    assign data[413]    =   { pl[1545],     pl[1546],   pl[1547],   pl[1548]    };
    assign data[414]    =   { pl[1549],     pl[1550],   pl[1551],   pl[1552]    };
    assign data[415]    =   { pl[1553],     pl[1554],   pl[1555],   pl[1556]    };
    assign data[416]    =   { pl[1557],     pl[1558],   pl[1559],   pl[1560]    };
    assign data[417]    =   { pl[1561],     pl[1562],   pl[1563],   pl[1564]    };
    assign data[418]    =   { pl[1565],     pl[1566],   pl[1567],   pl[1568]    };
    assign data[419]    =   { pl[1569],     pl[1570],   pl[1571],   pl[1572]    };
    assign data[420]    =   { pl[1573],     pl[1574],   pl[1575],   pl[1576]    };
    assign data[421]    =   { pl[1577],     pl[1578],   pl[1579],   pl[1580]    };
    assign data[422]    =   { pl[1581],     pl[1582],   pl[1583],   pl[1584]    };
    assign data[423]    =   { pl[1585],     pl[1586],   pl[1587],   pl[1588]    };
    assign data[424]    =   { pl[1589],     pl[1590],   pl[1591],   pl[1592]    };
    assign data[425]    =   { pl[1593],     pl[1594],   pl[1595],   pl[1596]    };
    assign data[426]    =   { pl[1597],     pl[1598],   pl[1599],   pl[1600]    };
    assign data[427]    =   { pl[1601],     pl[1602],   pl[1603],   pl[1604]    };
    assign data[428]    =   { pl[1605],     pl[1606],   pl[1607],   pl[1608]    };
    assign data[429]    =   { pl[1609],     pl[1610],   pl[1611],   pl[1612]    };
    assign data[430]    =   { pl[1613],     pl[1614],   pl[1615],   pl[1616]    };
    assign data[431]    =   { pl[1617],     pl[1618],   pl[1619],   pl[1620]    };
    assign data[432]    =   { pl[1621],     pl[1622],   pl[1623],   pl[1624]    };
    assign data[433]    =   { pl[1625],     pl[1626],   pl[1627],   pl[1628]    };
    assign data[434]    =   { pl[1629],     pl[1630],   pl[1631],   pl[1632]    };
    assign data[435]    =   { pl[1633],     pl[1634],   pl[1635],   pl[1636]    };
    assign data[436]    =   { pl[1637],     pl[1638],   pl[1639],   pl[1640]    };
    assign data[437]    =   { pl[1641],     pl[1642],   pl[1643],   pl[1644]    };
    assign data[438]    =   { pl[1645],     pl[1646],   pl[1647],   pl[1648]    };
    assign data[439]    =   { pl[1649],     pl[1650],   pl[1651],   pl[1652]    };
    assign data[440]    =   { pl[1653],     pl[1654],   pl[1655],   pl[1656]    };
    assign data[441]    =   { pl[1657],     pl[1658],   pl[1659],   pl[1660]    };
    assign data[442]    =   { pl[1661],     pl[1662],   pl[1663],   pl[1664]    };
    assign data[443]    =   { pl[1665],     pl[1666],   pl[1667],   pl[1668]    };
    assign data[444]    =   { pl[1669],     pl[1670],   pl[1671],   pl[1672]    };
    assign data[445]    =   { pl[1673],     pl[1674],   pl[1675],   pl[1676]    };
    assign data[446]    =   { pl[1677],     pl[1678],   pl[1679],   pl[1680]    };
    assign data[447]    =   { pl[1681],     pl[1682],   pl[1683],   pl[1684]    };
    assign data[448]    =   { pl[1685],     pl[1686],   pl[1687],   pl[1688]    };
    assign data[449]    =   { pl[1689],     pl[1690],   pl[1691],   pl[1692]    };
    assign data[450]    =   { pl[1693],     pl[1694],   pl[1695],   pl[1696]    };
    assign data[451]    =   { pl[1697],     pl[1698],   pl[1699],   pl[1700]    };
    assign data[452]    =   { pl[1701],     pl[1702],   pl[1703],   pl[1704]    };
    assign data[453]    =   { pl[1705],     pl[1706],   pl[1707],   pl[1708]    };
    assign data[454]    =   { pl[1709],     pl[1710],   pl[1711],   pl[1712]    };
    assign data[455]    =   { pl[1713],     pl[1714],   pl[1715],   pl[1716]    };
    assign data[456]    =   { pl[1717],     pl[1718],   pl[1719],   pl[1720]    };
    assign data[457]    =   { pl[1721],     pl[1722],   pl[1723],   pl[1724]    };
    assign data[458]    =   { pl[1725],     pl[1726],   pl[1727],   pl[1728]    };
    assign data[459]    =   { pl[1729],     pl[1730],   pl[1731],   pl[1732]    };
    assign data[460]    =   { pl[1733],     pl[1734],   pl[1735],   pl[1736]    };
    assign data[461]    =   { pl[1737],     pl[1738],   pl[1739],   pl[1740]    };
    assign data[462]    =   { pl[1741],     pl[1742],   pl[1743],   pl[1744]    };
    assign data[463]    =   { pl[1745],     pl[1746],   pl[1747],   pl[1748]    };
    assign data[464]    =   { pl[1749],     pl[1750],   pl[1751],   pl[1752]    };
    assign data[465]    =   { pl[1753],     pl[1754],   pl[1755],   pl[1756]    };
    assign data[466]    =   { pl[1757],     pl[1758],   pl[1759],   pl[1760]    };
    assign data[467]    =   { pl[1761],     pl[1762],   pl[1763],   pl[1764]    };
    assign data[468]    =   { pl[1765],     pl[1766],   pl[1767],   pl[1768]    };
    assign data[469]    =   { pl[1769],     pl[1770],   pl[1771],   pl[1772]    };
    assign data[470]    =   { pl[1773],     pl[1774],   pl[1775],   pl[1776]    };
    assign data[471]    =   { pl[1777],     pl[1778],   pl[1779],   pl[1780]    };
    assign data[472]    =   { pl[1781],     pl[1782],   pl[1783],   pl[1784]    };
    assign data[473]    =   { pl[1785],     pl[1786],   pl[1787],   pl[1788]    };
    assign data[474]    =   { pl[1789],     pl[1790],   pl[1791],   pl[1792]    };
    assign data[475]    =   { pl[1793],     pl[1794],   pl[1795],   pl[1796]    };
    assign data[476]    =   { pl[1797],     pl[1798],   pl[1799],   pl[1800]    };
    assign data[477]    =   { pl[1801],     pl[1802],   pl[1803],   pl[1804]    };
    assign data[478]    =   { pl[1805],     pl[1806],   pl[1807],   pl[1808]    };
    assign data[479]    =   { pl[1809],     pl[1810],   pl[1811],   pl[1812]    };
    assign data[480]    =   { pl[1813],     pl[1814],   pl[1815],   pl[1816]    };
    assign data[481]    =   { pl[1817],     pl[1818],   pl[1819],   pl[1820]    };
    assign data[482]    =   { pl[1821],     pl[1822],   pl[1823],   pl[1824]    };
    assign data[483]    =   { pl[1825],     pl[1826],   pl[1827],   pl[1828]    };
    assign data[484]    =   { pl[1829],     pl[1830],   pl[1831],   pl[1832]    };
    assign data[485]    =   { pl[1833],     pl[1834],   pl[1835],   pl[1836]    };
    assign data[486]    =   { pl[1837],     pl[1838],   pl[1839],   pl[1840]    };
    assign data[487]    =   { pl[1841],     pl[1842],   pl[1843],   pl[1844]    };
    assign data[488]    =   { pl[1845],     pl[1846],   pl[1847],   pl[1848]    };
    assign data[489]    =   { pl[1849],     pl[1850],   pl[1851],   pl[1852]    };
    assign data[490]    =   { pl[1853],     pl[1854],   pl[1855],   pl[1856]    };
    assign data[491]    =   { pl[1857],     pl[1858],   pl[1859],   pl[1860]    };
    assign data[492]    =   { pl[1861],     pl[1862],   pl[1863],   pl[1864]    };
    assign data[493]    =   { pl[1865],     pl[1866],   pl[1867],   pl[1868]    };
    assign data[494]    =   { pl[1869],     pl[1870],   pl[1871],   pl[1872]    };
    assign data[495]    =   { pl[1873],     pl[1874],   pl[1875],   pl[1876]    };
    assign data[496]    =   { pl[1877],     pl[1878],   pl[1879],   pl[1880]    };
    assign data[497]    =   { pl[1881],     pl[1882],   pl[1883],   pl[1884]    };
    assign data[498]    =   { pl[1885],     pl[1886],   pl[1887],   pl[1888]    };
    assign data[499]    =   { pl[1889],     pl[1890],   pl[1891],   pl[1892]    };
    assign data[500]    =   { pl[1893],     pl[1894],   pl[1895],   pl[1896]    };
    assign data[501]    =   { pl[1897],     pl[1898],   pl[1899],   fs[3]       };
    assign data[502]    =   { fec[96],      fec[97],    fec[98],    fec[99]     };
    assign data[503]    =   { fec[100],     fec[101],   fec[102],   fec[103]    };
    assign data[504]    =   { fec[104],     fec[105],   fec[106],   fec[107]    };
    assign data[505]    =   { fec[108],     fec[109],   fec[110],   fec[111]    };
    assign data[506]    =   { fec[112],     fec[113],   fec[114],   fec[115]    };
    assign data[507]    =   { fec[116],     fec[117],   fec[118],   fec[119]    };
    assign data[508]    =   { fec[120],     fec[121],   fec[122],   fec[123]    };
    assign data[509]    =   { fec[124],     fec[125],   fec[126],   fec[127]    };
    assign o_data   = data[i_address] ;

endmodule