`timescale 1 ns / 1 ps
//
// Copyright (c) 2016 by IP Cores, Inc.   All rights reserved.  This text
// contains proprietary, confidential information of IP Cores, Inc.,  and
// may be used, copied,  and/or disclosed only pursuant to the terms of a
// valid license agreement with IP Cores, Inc. This copyright notice must
// be retained as part of this text at all times.
//
// Rev. 1.0
//

module Kgmp16x128(
   input        [15:0] x,
   input       [127:0] y,
   output wire [127:0] z
);

   wire [7:0] Xo;
   wire [7:0] Xe;
   wire [63:0] Yo;
   wire [63:0] Ye;
   wire [71:0] Zo;
   wire [71:0] Ze;
   wire [71:0] Zeo;
   wire [71:0] z0;
   wire [71:0] z1;

   assign Xo = odd16(x);
   assign Xe = even16(x);

   assign Yo = odd128(y);
   assign Ye = even128(y);

   assign z0 = Ze ^ (Zo >> 1);
   assign z1 = Zeo ^ Ze ^ Zo;

   assign z = P128({48'h0, comb144( z0, z1)});

   Kgmp8x64 Pe (
      .x     ( Xe     ),
      .y     ( Ye     ),
      .z     ( Ze     )
   );

   Kgmp8x64 Po (
      .x     ( Xo     ),
      .y     ( Yo     ),
      .z     ( Zo     )
   );

   Kgmp8x64 Peo (
      .x     ( Xo ^ Xe   ),
      .y     ( Yo ^ Ye   ),
      .z     ( Zeo       )
   );

   function [63:0] odd128 (input [127:0] a);
      odd128 = { 
                 a[126], a[124], a[122], a[120], a[118], a[116], a[114], a[112], a[110], a[108], a[106], a[104], a[102], a[100], a[98], a[96],
                 a[94], a[92], a[90], a[88], a[86], a[84], a[82], a[80], a[78], a[76], a[74], a[72], a[70], a[68], a[66], a[64],
                 a[62], a[60], a[58], a[56], a[54], a[52], a[50], a[48], a[46], a[44], a[42], a[40], a[38], a[36], a[34], a[32],
                 a[30], a[28], a[26], a[24], a[22], a[20], a[18], a[16], a[14], a[12], a[10], a[8], a[6], a[4], a[2], a[0]
               };
   endfunction

   function [63:0] even128 (input [127:0] a);
      even128 = { 
                 a[127], a[125], a[123], a[121], a[119], a[117], a[115], a[113], a[111], a[109], a[107], a[105], a[103], a[101], a[99], a[97],
                 a[95], a[93], a[91], a[89], a[87], a[85], a[83], a[81], a[79], a[77], a[75], a[73], a[71], a[69], a[67], a[65],
                 a[63], a[61], a[59], a[57], a[55], a[53], a[51], a[49], a[47], a[45], a[43], a[41], a[39], a[37], a[35], a[33],
                 a[31], a[29], a[27], a[25], a[23], a[21], a[19], a[17], a[15], a[13], a[11], a[9], a[7], a[5], a[3], a[1]
                };
   endfunction

   function [7:0] odd16 (input [15:0] a);
      odd16  = { 
                 a[14], a[12], a[10], a[8], a[6], a[4], a[2], a[0]
               };
   endfunction

   function [7:0] even16 (input [15:0] a);
      even16  = {
                 a[15], a[13], a[11], a[9], a[7], a[5], a[3], a[1]
                };
   endfunction


   function [143:0] comb144 ( input [71:0] z0, input [71:0] z1 );
      comb144  = {
                   z0[71], z1[71], z0[70], z1[70], z0[69], z1[69], z0[68], z1[68],
                   z0[67], z1[67], z0[66], z1[66], z0[65], z1[65], z0[64], z1[64],
                   z0[63], z1[63], z0[62], z1[62], z0[61], z1[61], z0[60], z1[60],
                   z0[59], z1[59], z0[58], z1[58], z0[57], z1[57], z0[56], z1[56],
                   z0[55], z1[55], z0[54], z1[54], z0[53], z1[53], z0[52], z1[52],
                   z0[51], z1[51], z0[50], z1[50], z0[49], z1[49], z0[48], z1[48],
                   z0[47], z1[47], z0[46], z1[46], z0[45], z1[45], z0[44], z1[44],
                   z0[43], z1[43], z0[42], z1[42], z0[41], z1[41], z0[40], z1[40],
                   z0[39], z1[39], z0[38], z1[38], z0[37], z1[37], z0[36], z1[36],
                   z0[35], z1[35], z0[34], z1[34], z0[33], z1[33], z0[32], z1[32],
                   z0[31], z1[31], z0[30], z1[30], z0[29], z1[29], z0[28], z1[28],
                   z0[27], z1[27], z0[26], z1[26], z0[25], z1[25], z0[24], z1[24],
                   z0[23], z1[23], z0[22], z1[22], z0[21], z1[21], z0[20], z1[20],
                   z0[19], z1[19], z0[18], z1[18], z0[17], z1[17], z0[16], z1[16],
                   z0[15], z1[15], z0[14], z1[14], z0[13], z1[13], z0[12], z1[12],
                   z0[11], z1[11], z0[10], z1[10], z0[ 9], z1[ 9], z0[ 8], z1[ 8],
                   z0[ 7], z1[ 7], z0[ 6], z1[ 6], z0[ 5], z1[ 5], z0[ 4], z1[ 4],
                   z0[ 3], z1[ 3], z0[ 2], z1[ 2], z0[ 1], z1[ 1], z0[ 0], z1[ 0]
                };
   endfunction

// function [127:0] P128 (input [143:0] a);
//    P128 = {
//             a[63],
//             a[63] ^ a[62],
//             a[63] ^ a[62] ^ a[61],
//             a[62] ^ a[61] ^ a[60],
//             a[61] ^ a[60] ^ a[59],
//             a[60] ^ a[59] ^ a[58],
//             a[59] ^ a[58] ^ a[57],
//             a[63] ^ a[58] ^ a[57] ^ a[56],
//             a[62] ^ a[57] ^ a[56] ^ a[55],
//             a[61] ^ a[56] ^ a[55] ^ a[54],
//             a[60] ^ a[55] ^ a[54] ^ a[53],
//             a[59] ^ a[54] ^ a[53] ^ a[52],
//             a[58] ^ a[53] ^ a[52] ^ a[51],
//             a[57] ^ a[52] ^ a[51] ^ a[50],
//             a[56] ^ a[51] ^ a[50] ^ a[49],
//             a[55] ^ a[50] ^ a[49] ^ a[48],
//             a[54] ^ a[49] ^ a[48] ^ a[47],
//             a[53] ^ a[48] ^ a[47] ^ a[46],
//             a[52] ^ a[47] ^ a[46] ^ a[45],
//             a[51] ^ a[46] ^ a[45] ^ a[44],
//             a[50] ^ a[45] ^ a[44] ^ a[43],
//             a[49] ^ a[44] ^ a[43] ^ a[42],
//             a[48] ^ a[43] ^ a[42] ^ a[41],
//             a[47] ^ a[42] ^ a[41] ^ a[40],
//             a[46] ^ a[41] ^ a[40] ^ a[39],
//             a[45] ^ a[40] ^ a[39] ^ a[38],
//             a[44] ^ a[39] ^ a[38] ^ a[37],
//             a[43] ^ a[38] ^ a[37] ^ a[36],
//             a[42] ^ a[37] ^ a[36] ^ a[35],
//             a[41] ^ a[36] ^ a[35] ^ a[34],
//             a[40] ^ a[35] ^ a[34] ^ a[33],
//             a[39] ^ a[34] ^ a[33] ^ a[32],
//             a[38] ^ a[33] ^ a[32] ^ a[31],
//             a[37] ^ a[32] ^ a[31] ^ a[30],
//             a[36] ^ a[31] ^ a[30] ^ a[29],
//             a[35] ^ a[30] ^ a[29] ^ a[28],
//             a[34] ^ a[29] ^ a[28] ^ a[27],
//             a[33] ^ a[28] ^ a[27] ^ a[26],
//             a[32] ^ a[27] ^ a[26] ^ a[25],
//             a[31] ^ a[26] ^ a[25] ^ a[24],
//             a[30] ^ a[25] ^ a[24] ^ a[23],
//             a[29] ^ a[24] ^ a[23] ^ a[22],
//             a[28] ^ a[23] ^ a[22] ^ a[21],
//             a[27] ^ a[22] ^ a[21] ^ a[20],
//             a[26] ^ a[21] ^ a[20] ^ a[19],
//             a[25] ^ a[20] ^ a[19] ^ a[18],
//             a[24] ^ a[19] ^ a[18] ^ a[17],
//             a[23] ^ a[18] ^ a[17] ^ a[16],
//             a[143] ^ a[22] ^ a[17] ^ a[16] ^ a[15],
//             a[142] ^ a[21] ^ a[16] ^ a[15] ^ a[14],
//             a[141] ^ a[20] ^ a[15] ^ a[14] ^ a[13],
//             a[140] ^ a[19] ^ a[14] ^ a[13] ^ a[12],
//             a[139] ^ a[18] ^ a[13] ^ a[12] ^ a[11],
//             a[138] ^ a[17] ^ a[12] ^ a[11] ^ a[10],
//             a[137] ^ a[16] ^ a[11] ^ a[10] ^ a[9],
//             a[136] ^ a[15] ^ a[10] ^ a[9] ^ a[8],
//             a[135] ^ a[14] ^ a[9] ^ a[8] ^ a[7],
//             a[134] ^ a[13] ^ a[8] ^ a[7] ^ a[6],
//             a[133] ^ a[12] ^ a[7] ^ a[6] ^ a[5],
//             a[132] ^ a[11] ^ a[6] ^ a[5] ^ a[4],
//             a[131] ^ a[10] ^ a[5] ^ a[4] ^ a[3],
//             a[130] ^ a[9] ^ a[4] ^ a[3] ^ a[2],
//             a[129] ^ a[8] ^ a[3] ^ a[2] ^ a[1],
//             a[128] ^ a[7] ^ a[2] ^ a[1] ^ a[0],
//             a[127] ^ a[6] ^ a[1] ^ a[0],
//             a[126] ^ a[5] ^ a[0],
//             a[125] ^ a[4],
//             a[124] ^ a[3],
//             a[123] ^ a[2],
//             a[122] ^ a[1],
//             a[121] ^ a[0],
//             a[120:64]
//           };
// endfunction

   function [127:0] P128 (input [143:0] a);
      P128 = {
                   a[143] ^ a[15],
                   a[142] ^ a[15] ^ a[14],
                   a[141] ^ a[15] ^ a[14] ^ a[13],
                   a[140] ^ a[14] ^ a[13] ^ a[12],
                   a[139] ^ a[13] ^ a[12] ^ a[11],
                   a[138] ^ a[12] ^ a[11] ^ a[10],
                   a[137] ^ a[11] ^ a[10] ^ a[9],
                   a[136] ^ a[15] ^ a[10] ^ a[9] ^ a[8],
                   a[135] ^ a[14] ^ a[9] ^ a[8] ^ a[7],
                   a[134] ^ a[13] ^ a[8] ^ a[7] ^ a[6],
                   a[133] ^ a[12] ^ a[7] ^ a[6] ^ a[5],
                   a[132] ^ a[11] ^ a[6] ^ a[5] ^ a[4],
                   a[131] ^ a[10] ^ a[5] ^ a[4] ^ a[3],
                   a[130] ^ a[9] ^ a[4] ^ a[3] ^ a[2],
                   a[129] ^ a[8] ^ a[3] ^ a[2] ^ a[1],
                   a[128] ^ a[7] ^ a[2] ^ a[1] ^ a[0],
                   a[127] ^ a[6] ^ a[1] ^ a[0],
                   a[126] ^ a[5] ^ a[0],
                   a[125] ^ a[4],
                   a[124] ^ a[3],
                   a[123] ^ a[2],
                   a[122] ^ a[1],
                   a[121] ^ a[0],
                   a[120:16]
             };
   endfunction


endmodule
