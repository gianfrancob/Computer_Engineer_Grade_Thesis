module tb_autogen_gcm_aes
(
    // OUTPUTS.
    output      wire                    o_compOK                                            ,
    output      wire                    o_ciphertextOK                                      ,
    output      wire                    o_tagOK
    // INPUTS.
    // none so far
);

// LOCALPARAMETERS.
// ----------------------------------------------------------------------------------------------------
localparam                              NB_BLOCK                =   128                     ;
localparam                              N_BLOCKS                =   2                       ;
localparam                              NB_DATA                 =   N_BLOCKS*NB_BLOCK       ;
localparam                              NB_IV                   =   96                      ;
localparam                              NB_KEY                  =   256                     ;
localparam                              NB_INC_MODE             =   2                       ;
localparam                              USE_LUT_IN_SUBBYTES     =   0                       ;
localparam                              NB_N_MESSAGES           =   10                      ;
localparam                              RUN_TIME                =   1240                      ;


// INTERNAL SIGNALS.
// ----------------------------------------------------------------------------------------------------
wire                                    tb_i_valid                      [ RUN_TIME-1:0  ]   ;
wire                                    tb_i_reset                      [ RUN_TIME-1:0  ]   ;
wire                                    tb_i_sop                        [ RUN_TIME-1:0  ]   ;
wire                                    tb_i_key_update                 [ RUN_TIME-1:0  ]   ;
wire    [ NB_KEY-1:0        ]           tb_i_key                        [ RUN_TIME-1:0  ]   ;
wire    [ NB_IV-1:0         ]           tb_i_iv                         [ RUN_TIME-1:0  ]   ;
wire    [ NB_BLOCK/2-1:0    ]           tb_i_rf_static_aad_length       [ RUN_TIME-1:0  ]   ;
wire    [ NB_DATA-1:0       ]           tb_i_aad                        [ RUN_TIME-1:0  ]   ;
wire    [ NB_BLOCK/2-1:0    ]           tb_i_rf_static_plaintext_length [ RUN_TIME-1:0  ]   ;
wire    [ NB_DATA-1:0       ]           tb_i_plaintext                  [ RUN_TIME-1:0  ]   ;
wire    [ NB_INC_MODE-1:0   ]           tb_i_rf_static_inc_mode                             ;
wire                                    tb_i_rf_mode_gmac               [ RUN_TIME-1:0  ]   ;
wire                                    tb_i_rf_static_encrypt          [ RUN_TIME-1:0  ]   ;
wire                                    tb_i_clear_fault_flags          [ RUN_TIME-1:0  ]   ;
wire    [ NB_DATA-1:0       ]           tb_o_ciphertext                 [ RUN_TIME-1:0  ]   ;
wire                                    tb_o_fail                       [ RUN_TIME-1:0  ]   ;
wire                                    tb_o_sop                        [ RUN_TIME-1:0  ]   ;
wire                                    tb_o_valid                      [ RUN_TIME-1:0  ]   ;
wire    [ NB_BLOCK-1:0      ]           tb_o_tag                        [ RUN_TIME-1:0  ]   ;
wire                                    tb_o_tag_ready                  [ RUN_TIME-1:0  ]   ;

wire    [ NB_DATA-1:0       ]           tb_gcm_aes_core_o_ciphertext                        ;
wire                                    tb_gcm_aes_core_o_fail                              ;
wire                                    tb_gcm_aes_core_o_sop                               ;
wire                                    tb_gcm_aes_core_o_valid                             ;
wire    [ NB_BLOCK-1:0      ]           tb_gcm_aes_core_o_tag                               ;
wire                                    tb_gcm_aes_core_o_tag_ready                         ;
wire                                    tb_gcm_aes_core_o_fault_sop_and_keyupdate           ;

reg                                     tb_i_clock                                          ;

wire    [ NB_DATA-1:0       ]           o_ciphertext                                        ;
wire                                    o_sop                                               ;
wire                                    o_valid                                             ;
wire    [ NB_BLOCK-1:0      ]           o_tag                                               ;
wire                                    o_tag_ready                                         ;
wire    [ NB_KEY-1:0        ]           i_key                                               ;
wire    [ NB_DATA-1:0       ]           i_plaintext                                         ;
wire    [ NB_DATA-1:0       ]           i_aad                                               ;
wire    [ NB_IV-1:0         ]           i_iv                                                ;
wire    [ NB_BLOCK/2-1:0    ]           i_rf_static_aad_length                              ;
wire    [ NB_BLOCK/2-1:0    ]           i_rf_static_plaintext_length                        ;
wire                                    i_sop                                               ;
wire                                    i_valid                                             ;
wire                                    i_key_update                                        ;
wire                                    i_rf_mode_gmac                                      ;
wire                                    i_rf_static_encrypt                                 ;
wire                                    i_clear_fault_flags                                 ;
wire                                    i_reset                                             ;

reg                                     o_ciphertextOK_reg                                  ;
reg                                     o_tagOK_reg                                         ;

integer                                 clock_ctr                                           ;


// MISC.
// ----------------------------------------------------------------------------------------------------
initial begin
    tb_i_clock  <= 0    ;
    clock_ctr   <= 0    ;
end

always #5 tb_i_clock    <= ~tb_i_clock  ;

always @( posedge tb_i_clock )
begin
    clock_ctr   <= clock_ctr + 1    ;
    if ( clock_ctr == RUN_TIME + 1 )
        $stop();
end

assign  o_ciphertext                    = tb_o_ciphertext                   [clock_ctr] ;
assign  o_sop                           = tb_o_sop                          [clock_ctr] ;
assign  o_valid                         = tb_o_valid                        [clock_ctr] ;
assign  o_tag                           = tb_o_tag                          [clock_ctr] ;
assign  o_tag_ready                     = tb_o_tag_ready                    [clock_ctr] ;
assign  tb_i_rf_static_inc_mode         = 2'd2                                          ;
assign  i_plaintext                     = tb_i_plaintext                    [clock_ctr] ;
assign  i_key                           = tb_i_key                          [clock_ctr] ;
assign  i_aad                           = tb_i_aad                          [clock_ctr] ;
assign  i_iv                            = tb_i_iv                           [clock_ctr] ;
assign  i_rf_static_aad_length          = tb_i_rf_static_aad_length         [clock_ctr] ;
assign  i_rf_static_plaintext_length    = tb_i_rf_static_plaintext_length   [clock_ctr] ;
assign  i_sop                           = tb_i_sop                          [clock_ctr] ;
assign  i_valid                         = tb_i_valid                        [clock_ctr] ;
assign  i_key_update                    = tb_i_key_update                   [clock_ctr] ;
assign  i_rf_mode_gmac                  = tb_i_rf_mode_gmac                 [clock_ctr] ;
assign  i_rf_static_encrypt             = tb_i_rf_static_encrypt            [clock_ctr] ;
assign  i_clear_fault_flags             = tb_i_clear_fault_flags            [clock_ctr] ;
assign  i_reset                         = tb_i_reset                        [clock_ctr] ;


// COMPS.
// ----------------------------------------------------------------------------------------------------
always @( posedge tb_i_clock )
begin
    if (o_valid)
        if (i_rf_static_plaintext_length[7])
            o_ciphertextOK_reg  <=  (tb_gcm_aes_core_o_ciphertext[0+:128] == o_ciphertext[0+:128])  ;
        else
            o_ciphertextOK_reg  <=  (tb_gcm_aes_core_o_ciphertext == o_ciphertext)  ;
end

assign  o_ciphertextOK  =   (tb_gcm_aes_core_o_valid)   ?
                            ( (i_rf_static_plaintext_length[7])   ?
                            (tb_gcm_aes_core_o_ciphertext[0+:128] == o_ciphertext[0+:128]) :
                            (tb_gcm_aes_core_o_ciphertext == o_ciphertext) ) : o_ciphertextOK_reg   ;

always @( posedge tb_i_clock )
begin
    if (o_tag_ready)
        o_tagOK_reg     <=  (tb_gcm_aes_core_o_tag == o_tag)    ;
end

assign  o_tagOK         =   (tb_gcm_aes_core_o_tag_ready)   ?
                            (tb_gcm_aes_core_o_tag == o_tag) : o_tagOK_reg  ;

assign  o_compOK        =   (o_ciphertextOK == 1'b1) & (o_tagOK == 1'b1)    ;


// GCM AES CORE.
// ----------------------------------------------------------------------------------------------------
gcm_aes_core
#(
    .NB_BLOCK                       ( NB_BLOCK                                      ),
    .N_BLOCKS                       ( N_BLOCKS                                      ),
    .NB_DATA                        ( NB_DATA                                       ),
    .NB_KEY                         ( NB_KEY                                        ),
    .NB_IV                          ( NB_IV                                         ),
    .NB_INC_MODE                    ( NB_INC_MODE                                   ),
    .USE_LUT_IN_SUBBYTES            ( USE_LUT_IN_SUBBYTES                           ),
    .NB_N_MESSAGES                  ( NB_N_MESSAGES                                 )
)
u_gcm_aes_core_cipher
(
    .o_ciphertext                   ( tb_gcm_aes_core_o_ciphertext                  ),
    .o_fail                         ( tb_gcm_aes_core_o_fail                        ),
    .o_sop                          ( tb_gcm_aes_core_o_sop                         ),
    .o_valid                        ( tb_gcm_aes_core_o_valid                       ),
    .o_tag                          ( tb_gcm_aes_core_o_tag                         ),
    .o_tag_ready                    ( tb_gcm_aes_core_o_tag_ready                   ),
    .o_fault_sop_and_keyupdate      ( tb_gcm_aes_core_o_fault_sop_and_keyupdate     ),
    .i_plaintext                    ( i_plaintext                                   ),
    .i_tag                          ( /*unused*/                                    ),
    .i_tag_ready                    ( /*unused*/                                    ),
    .i_rf_static_key                ( i_key                                         ),
    .i_rf_static_aad                ( i_aad                                         ),
    .i_rf_static_iv                 ( i_iv                                          ),
    .i_rf_static_length_aad         ( i_rf_static_aad_length                        ),
    .i_rf_static_length_plaintext   ( i_rf_static_plaintext_length                  ),
    .i_sop                          ( i_sop                                         ),
    .i_valid                        ( i_valid                                       ),
    .i_enable                       ( 1'b1                                          ),
    .i_update_key                   ( i_key_update                                  ),
    .i_rf_static_inc_mode           ( tb_i_rf_static_inc_mode                       ),
    .i_rf_mode_gmac                 ( i_rf_mode_gmac                                ),
    .i_rf_static_encrypt            ( i_rf_static_encrypt                           ),
    .i_clear_fault_flags            ( i_clear_fault_flags                           ),
    .i_reset                        ( i_reset                                       ),
    .i_clock                        ( tb_i_clock                                    )
);


// AUTOGENERATED VECTORS.
// ----------------------------------------------------------------------------------------------------
// CLK no. 0/1240
// *************************************************
assign   tb_i_valid[0]                      =   1'b0;
assign   tb_i_reset[0]                      =   1'b1;
assign   tb_i_sop[0]                        =   1'b0;
assign   tb_i_key_update[0]                 =   1'b0;
assign   tb_i_key[0]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[0]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[0]               =   1'b0;
assign   tb_i_rf_static_encrypt[0]          =   1'b1;
assign   tb_i_clear_fault_flags[0]          =   1'b0;
assign   tb_i_rf_static_aad_length[0]       =   64'h0000000000000100;
assign   tb_i_aad[0]                        =   tb_i_aad[0];
assign   tb_i_rf_static_plaintext_length[0] =   64'h0000000000000200;
assign   tb_i_plaintext[0]                  =   tb_i_plaintext[0];
assign   tb_o_valid[0]                      =   1'b0;
assign   tb_o_sop[0]                        =   1'b0;
assign   tb_o_ciphertext[0]                 =   tb_o_ciphertext[0];
assign   tb_o_tag_ready[0]                  =   1'b0;
assign   tb_o_tag[0]                        =   tb_o_tag[0];

// CLK no. 1/1240
// *************************************************
assign   tb_i_valid[1]                      =   1'b0;
assign   tb_i_reset[1]                      =   1'b0;
assign   tb_i_sop[1]                        =   1'b1;
assign   tb_i_key_update[1]                 =   1'b1;
assign   tb_i_key[1]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1]               =   1'b0;
assign   tb_i_rf_static_encrypt[1]          =   1'b1;
assign   tb_i_clear_fault_flags[1]          =   1'b0;
assign   tb_i_rf_static_aad_length[1]       =   64'h0000000000000100;
assign   tb_i_aad[1]                        =   tb_i_aad[0];
assign   tb_i_rf_static_plaintext_length[1] =   64'h0000000000000200;
assign   tb_i_plaintext[1]                  =   tb_i_plaintext[0];
assign   tb_o_valid[1]                      =   1'b0;
assign   tb_o_sop[1]                        =   1'b0;
assign   tb_o_ciphertext[1]                 =   tb_o_ciphertext[0];
assign   tb_o_tag_ready[1]                  =   1'b0;
assign   tb_o_tag[1]                        =   tb_o_tag[0];

// CLK no. 2/1240
// *************************************************
assign   tb_i_valid[2]                      =   1'b1;
assign   tb_i_reset[2]                      =   1'b0;
assign   tb_i_sop[2]                        =   1'b0;
assign   tb_i_key_update[2]                 =   1'b0;
assign   tb_i_key[2]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[2]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[2]               =   1'b0;
assign   tb_i_rf_static_encrypt[2]          =   1'b1;
assign   tb_i_clear_fault_flags[2]          =   1'b0;
assign   tb_i_rf_static_aad_length[2]       =   64'h0000000000000100;
assign   tb_i_aad[2]                        =   256'h5999366a10a3ca7ab06bc4cb4b64d7e68db6b469c41d0619b4ff00b0ed2a2ae3;
assign   tb_i_rf_static_plaintext_length[2] =   64'h0000000000000200;
assign   tb_i_plaintext[2]                  =   tb_i_plaintext[1];
assign   tb_o_valid[2]                      =   1'b0;
assign   tb_o_sop[2]                        =   1'b0;
assign   tb_o_ciphertext[2]                 =   tb_o_ciphertext[1];
assign   tb_o_tag_ready[2]                  =   1'b0;
assign   tb_o_tag[2]                        =   tb_o_tag[1];

// CLK no. 3/1240
// *************************************************
assign   tb_i_valid[3]                      =   1'b1;
assign   tb_i_reset[3]                      =   1'b0;
assign   tb_i_sop[3]                        =   1'b0;
assign   tb_i_key_update[3]                 =   1'b0;
assign   tb_i_key[3]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[3]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[3]               =   1'b0;
assign   tb_i_rf_static_encrypt[3]          =   1'b1;
assign   tb_i_clear_fault_flags[3]          =   1'b0;
assign   tb_i_rf_static_aad_length[3]       =   64'h0000000000000100;
assign   tb_i_aad[3]                        =   tb_i_aad[2];
assign   tb_i_rf_static_plaintext_length[3] =   64'h0000000000000200;
assign   tb_i_plaintext[3]                  =   256'hbf83800a673ca6524f6147781ecf858a03dd13090e7476ab712349d2c51fe3dc;
assign   tb_o_valid[3]                      =   1'b0;
assign   tb_o_sop[3]                        =   1'b0;
assign   tb_o_ciphertext[3]                 =   tb_o_ciphertext[2];
assign   tb_o_tag_ready[3]                  =   1'b0;
assign   tb_o_tag[3]                        =   tb_o_tag[2];

// CLK no. 4/1240
// *************************************************
assign   tb_i_valid[4]                      =   1'b1;
assign   tb_i_reset[4]                      =   1'b0;
assign   tb_i_sop[4]                        =   1'b0;
assign   tb_i_key_update[4]                 =   1'b0;
assign   tb_i_key[4]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[4]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[4]               =   1'b0;
assign   tb_i_rf_static_encrypt[4]          =   1'b1;
assign   tb_i_clear_fault_flags[4]          =   1'b0;
assign   tb_i_rf_static_aad_length[4]       =   64'h0000000000000100;
assign   tb_i_aad[4]                        =   tb_i_aad[3];
assign   tb_i_rf_static_plaintext_length[4] =   64'h0000000000000200;
assign   tb_i_plaintext[4]                  =   256'h09653965c6cb10294b8ea6e0948f4f3cff4c2b629311a5e04fdc9279111fcd88;
assign   tb_o_valid[4]                      =   1'b0;
assign   tb_o_sop[4]                        =   1'b0;
assign   tb_o_ciphertext[4]                 =   tb_o_ciphertext[3];
assign   tb_o_tag_ready[4]                  =   1'b0;
assign   tb_o_tag[4]                        =   tb_o_tag[3];

// CLK no. 5/1240
// *************************************************
assign   tb_i_valid[5]                      =   1'b0;
assign   tb_i_reset[5]                      =   1'b0;
assign   tb_i_sop[5]                        =   1'b0;
assign   tb_i_key_update[5]                 =   1'b0;
assign   tb_i_key[5]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[5]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[5]               =   1'b0;
assign   tb_i_rf_static_encrypt[5]          =   1'b1;
assign   tb_i_clear_fault_flags[5]          =   1'b0;
assign   tb_i_rf_static_aad_length[5]       =   64'h0000000000000100;
assign   tb_i_aad[5]                        =   tb_i_aad[4];
assign   tb_i_rf_static_plaintext_length[5] =   64'h0000000000000200;
assign   tb_i_plaintext[5]                  =   tb_i_plaintext[4];
assign   tb_o_valid[5]                      =   1'b0;
assign   tb_o_sop[5]                        =   1'b0;
assign   tb_o_ciphertext[5]                 =   tb_o_ciphertext[4];
assign   tb_o_tag_ready[5]                  =   1'b0;
assign   tb_o_tag[5]                        =   tb_o_tag[4];

// CLK no. 6/1240
// *************************************************
assign   tb_i_valid[6]                      =   1'b0;
assign   tb_i_reset[6]                      =   1'b0;
assign   tb_i_sop[6]                        =   1'b0;
assign   tb_i_key_update[6]                 =   1'b0;
assign   tb_i_key[6]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[6]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[6]               =   1'b0;
assign   tb_i_rf_static_encrypt[6]          =   1'b1;
assign   tb_i_clear_fault_flags[6]          =   1'b0;
assign   tb_i_rf_static_aad_length[6]       =   64'h0000000000000100;
assign   tb_i_aad[6]                        =   tb_i_aad[5];
assign   tb_i_rf_static_plaintext_length[6] =   64'h0000000000000200;
assign   tb_i_plaintext[6]                  =   tb_i_plaintext[5];
assign   tb_o_valid[6]                      =   1'b0;
assign   tb_o_sop[6]                        =   1'b0;
assign   tb_o_ciphertext[6]                 =   tb_o_ciphertext[5];
assign   tb_o_tag_ready[6]                  =   1'b0;
assign   tb_o_tag[6]                        =   tb_o_tag[5];

// CLK no. 7/1240
// *************************************************
assign   tb_i_valid[7]                      =   1'b0;
assign   tb_i_reset[7]                      =   1'b0;
assign   tb_i_sop[7]                        =   1'b0;
assign   tb_i_key_update[7]                 =   1'b0;
assign   tb_i_key[7]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[7]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[7]               =   1'b0;
assign   tb_i_rf_static_encrypt[7]          =   1'b1;
assign   tb_i_clear_fault_flags[7]          =   1'b0;
assign   tb_i_rf_static_aad_length[7]       =   64'h0000000000000100;
assign   tb_i_aad[7]                        =   tb_i_aad[6];
assign   tb_i_rf_static_plaintext_length[7] =   64'h0000000000000200;
assign   tb_i_plaintext[7]                  =   tb_i_plaintext[6];
assign   tb_o_valid[7]                      =   1'b0;
assign   tb_o_sop[7]                        =   1'b0;
assign   tb_o_ciphertext[7]                 =   tb_o_ciphertext[6];
assign   tb_o_tag_ready[7]                  =   1'b0;
assign   tb_o_tag[7]                        =   tb_o_tag[6];

// CLK no. 8/1240
// *************************************************
assign   tb_i_valid[8]                      =   1'b0;
assign   tb_i_reset[8]                      =   1'b0;
assign   tb_i_sop[8]                        =   1'b0;
assign   tb_i_key_update[8]                 =   1'b0;
assign   tb_i_key[8]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[8]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[8]               =   1'b0;
assign   tb_i_rf_static_encrypt[8]          =   1'b1;
assign   tb_i_clear_fault_flags[8]          =   1'b0;
assign   tb_i_rf_static_aad_length[8]       =   64'h0000000000000100;
assign   tb_i_aad[8]                        =   tb_i_aad[7];
assign   tb_i_rf_static_plaintext_length[8] =   64'h0000000000000200;
assign   tb_i_plaintext[8]                  =   tb_i_plaintext[7];
assign   tb_o_valid[8]                      =   1'b0;
assign   tb_o_sop[8]                        =   1'b0;
assign   tb_o_ciphertext[8]                 =   tb_o_ciphertext[7];
assign   tb_o_tag_ready[8]                  =   1'b0;
assign   tb_o_tag[8]                        =   tb_o_tag[7];

// CLK no. 9/1240
// *************************************************
assign   tb_i_valid[9]                      =   1'b0;
assign   tb_i_reset[9]                      =   1'b0;
assign   tb_i_sop[9]                        =   1'b0;
assign   tb_i_key_update[9]                 =   1'b0;
assign   tb_i_key[9]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[9]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[9]               =   1'b0;
assign   tb_i_rf_static_encrypt[9]          =   1'b1;
assign   tb_i_clear_fault_flags[9]          =   1'b0;
assign   tb_i_rf_static_aad_length[9]       =   64'h0000000000000100;
assign   tb_i_aad[9]                        =   tb_i_aad[8];
assign   tb_i_rf_static_plaintext_length[9] =   64'h0000000000000200;
assign   tb_i_plaintext[9]                  =   tb_i_plaintext[8];
assign   tb_o_valid[9]                      =   1'b0;
assign   tb_o_sop[9]                        =   1'b0;
assign   tb_o_ciphertext[9]                 =   tb_o_ciphertext[8];
assign   tb_o_tag_ready[9]                  =   1'b0;
assign   tb_o_tag[9]                        =   tb_o_tag[8];

// CLK no. 10/1240
// *************************************************
assign   tb_i_valid[10]                      =   1'b0;
assign   tb_i_reset[10]                      =   1'b0;
assign   tb_i_sop[10]                        =   1'b0;
assign   tb_i_key_update[10]                 =   1'b0;
assign   tb_i_key[10]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[10]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[10]               =   1'b0;
assign   tb_i_rf_static_encrypt[10]          =   1'b1;
assign   tb_i_clear_fault_flags[10]          =   1'b0;
assign   tb_i_rf_static_aad_length[10]       =   64'h0000000000000100;
assign   tb_i_aad[10]                        =   tb_i_aad[9];
assign   tb_i_rf_static_plaintext_length[10] =   64'h0000000000000200;
assign   tb_i_plaintext[10]                  =   tb_i_plaintext[9];
assign   tb_o_valid[10]                      =   1'b0;
assign   tb_o_sop[10]                        =   1'b0;
assign   tb_o_ciphertext[10]                 =   tb_o_ciphertext[9];
assign   tb_o_tag_ready[10]                  =   1'b0;
assign   tb_o_tag[10]                        =   tb_o_tag[9];

// CLK no. 11/1240
// *************************************************
assign   tb_i_valid[11]                      =   1'b0;
assign   tb_i_reset[11]                      =   1'b0;
assign   tb_i_sop[11]                        =   1'b0;
assign   tb_i_key_update[11]                 =   1'b0;
assign   tb_i_key[11]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[11]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[11]               =   1'b0;
assign   tb_i_rf_static_encrypt[11]          =   1'b1;
assign   tb_i_clear_fault_flags[11]          =   1'b0;
assign   tb_i_rf_static_aad_length[11]       =   64'h0000000000000100;
assign   tb_i_aad[11]                        =   tb_i_aad[10];
assign   tb_i_rf_static_plaintext_length[11] =   64'h0000000000000200;
assign   tb_i_plaintext[11]                  =   tb_i_plaintext[10];
assign   tb_o_valid[11]                      =   1'b0;
assign   tb_o_sop[11]                        =   1'b0;
assign   tb_o_ciphertext[11]                 =   tb_o_ciphertext[10];
assign   tb_o_tag_ready[11]                  =   1'b0;
assign   tb_o_tag[11]                        =   tb_o_tag[10];

// CLK no. 12/1240
// *************************************************
assign   tb_i_valid[12]                      =   1'b0;
assign   tb_i_reset[12]                      =   1'b0;
assign   tb_i_sop[12]                        =   1'b0;
assign   tb_i_key_update[12]                 =   1'b0;
assign   tb_i_key[12]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[12]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[12]               =   1'b0;
assign   tb_i_rf_static_encrypt[12]          =   1'b1;
assign   tb_i_clear_fault_flags[12]          =   1'b0;
assign   tb_i_rf_static_aad_length[12]       =   64'h0000000000000100;
assign   tb_i_aad[12]                        =   tb_i_aad[11];
assign   tb_i_rf_static_plaintext_length[12] =   64'h0000000000000200;
assign   tb_i_plaintext[12]                  =   tb_i_plaintext[11];
assign   tb_o_valid[12]                      =   1'b0;
assign   tb_o_sop[12]                        =   1'b0;
assign   tb_o_ciphertext[12]                 =   tb_o_ciphertext[11];
assign   tb_o_tag_ready[12]                  =   1'b0;
assign   tb_o_tag[12]                        =   tb_o_tag[11];

// CLK no. 13/1240
// *************************************************
assign   tb_i_valid[13]                      =   1'b0;
assign   tb_i_reset[13]                      =   1'b0;
assign   tb_i_sop[13]                        =   1'b0;
assign   tb_i_key_update[13]                 =   1'b0;
assign   tb_i_key[13]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[13]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[13]               =   1'b0;
assign   tb_i_rf_static_encrypt[13]          =   1'b1;
assign   tb_i_clear_fault_flags[13]          =   1'b0;
assign   tb_i_rf_static_aad_length[13]       =   64'h0000000000000100;
assign   tb_i_aad[13]                        =   tb_i_aad[12];
assign   tb_i_rf_static_plaintext_length[13] =   64'h0000000000000200;
assign   tb_i_plaintext[13]                  =   tb_i_plaintext[12];
assign   tb_o_valid[13]                      =   1'b0;
assign   tb_o_sop[13]                        =   1'b0;
assign   tb_o_ciphertext[13]                 =   tb_o_ciphertext[12];
assign   tb_o_tag_ready[13]                  =   1'b0;
assign   tb_o_tag[13]                        =   tb_o_tag[12];

// CLK no. 14/1240
// *************************************************
assign   tb_i_valid[14]                      =   1'b0;
assign   tb_i_reset[14]                      =   1'b0;
assign   tb_i_sop[14]                        =   1'b0;
assign   tb_i_key_update[14]                 =   1'b0;
assign   tb_i_key[14]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[14]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[14]               =   1'b0;
assign   tb_i_rf_static_encrypt[14]          =   1'b1;
assign   tb_i_clear_fault_flags[14]          =   1'b0;
assign   tb_i_rf_static_aad_length[14]       =   64'h0000000000000100;
assign   tb_i_aad[14]                        =   tb_i_aad[13];
assign   tb_i_rf_static_plaintext_length[14] =   64'h0000000000000200;
assign   tb_i_plaintext[14]                  =   tb_i_plaintext[13];
assign   tb_o_valid[14]                      =   1'b0;
assign   tb_o_sop[14]                        =   1'b0;
assign   tb_o_ciphertext[14]                 =   tb_o_ciphertext[13];
assign   tb_o_tag_ready[14]                  =   1'b0;
assign   tb_o_tag[14]                        =   tb_o_tag[13];

// CLK no. 15/1240
// *************************************************
assign   tb_i_valid[15]                      =   1'b0;
assign   tb_i_reset[15]                      =   1'b0;
assign   tb_i_sop[15]                        =   1'b0;
assign   tb_i_key_update[15]                 =   1'b0;
assign   tb_i_key[15]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[15]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[15]               =   1'b0;
assign   tb_i_rf_static_encrypt[15]          =   1'b1;
assign   tb_i_clear_fault_flags[15]          =   1'b0;
assign   tb_i_rf_static_aad_length[15]       =   64'h0000000000000100;
assign   tb_i_aad[15]                        =   tb_i_aad[14];
assign   tb_i_rf_static_plaintext_length[15] =   64'h0000000000000200;
assign   tb_i_plaintext[15]                  =   tb_i_plaintext[14];
assign   tb_o_valid[15]                      =   1'b0;
assign   tb_o_sop[15]                        =   1'b0;
assign   tb_o_ciphertext[15]                 =   tb_o_ciphertext[14];
assign   tb_o_tag_ready[15]                  =   1'b0;
assign   tb_o_tag[15]                        =   tb_o_tag[14];

// CLK no. 16/1240
// *************************************************
assign   tb_i_valid[16]                      =   1'b0;
assign   tb_i_reset[16]                      =   1'b0;
assign   tb_i_sop[16]                        =   1'b0;
assign   tb_i_key_update[16]                 =   1'b0;
assign   tb_i_key[16]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[16]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[16]               =   1'b0;
assign   tb_i_rf_static_encrypt[16]          =   1'b1;
assign   tb_i_clear_fault_flags[16]          =   1'b0;
assign   tb_i_rf_static_aad_length[16]       =   64'h0000000000000100;
assign   tb_i_aad[16]                        =   tb_i_aad[15];
assign   tb_i_rf_static_plaintext_length[16] =   64'h0000000000000200;
assign   tb_i_plaintext[16]                  =   tb_i_plaintext[15];
assign   tb_o_valid[16]                      =   1'b0;
assign   tb_o_sop[16]                        =   1'b0;
assign   tb_o_ciphertext[16]                 =   tb_o_ciphertext[15];
assign   tb_o_tag_ready[16]                  =   1'b0;
assign   tb_o_tag[16]                        =   tb_o_tag[15];

// CLK no. 17/1240
// *************************************************
assign   tb_i_valid[17]                      =   1'b0;
assign   tb_i_reset[17]                      =   1'b0;
assign   tb_i_sop[17]                        =   1'b0;
assign   tb_i_key_update[17]                 =   1'b0;
assign   tb_i_key[17]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[17]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[17]               =   1'b0;
assign   tb_i_rf_static_encrypt[17]          =   1'b1;
assign   tb_i_clear_fault_flags[17]          =   1'b0;
assign   tb_i_rf_static_aad_length[17]       =   64'h0000000000000100;
assign   tb_i_aad[17]                        =   tb_i_aad[16];
assign   tb_i_rf_static_plaintext_length[17] =   64'h0000000000000200;
assign   tb_i_plaintext[17]                  =   tb_i_plaintext[16];
assign   tb_o_valid[17]                      =   1'b0;
assign   tb_o_sop[17]                        =   1'b0;
assign   tb_o_ciphertext[17]                 =   tb_o_ciphertext[16];
assign   tb_o_tag_ready[17]                  =   1'b0;
assign   tb_o_tag[17]                        =   tb_o_tag[16];

// CLK no. 18/1240
// *************************************************
assign   tb_i_valid[18]                      =   1'b0;
assign   tb_i_reset[18]                      =   1'b0;
assign   tb_i_sop[18]                        =   1'b0;
assign   tb_i_key_update[18]                 =   1'b0;
assign   tb_i_key[18]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[18]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[18]               =   1'b0;
assign   tb_i_rf_static_encrypt[18]          =   1'b1;
assign   tb_i_clear_fault_flags[18]          =   1'b0;
assign   tb_i_rf_static_aad_length[18]       =   64'h0000000000000100;
assign   tb_i_aad[18]                        =   tb_i_aad[17];
assign   tb_i_rf_static_plaintext_length[18] =   64'h0000000000000200;
assign   tb_i_plaintext[18]                  =   tb_i_plaintext[17];
assign   tb_o_valid[18]                      =   1'b0;
assign   tb_o_sop[18]                        =   1'b0;
assign   tb_o_ciphertext[18]                 =   tb_o_ciphertext[17];
assign   tb_o_tag_ready[18]                  =   1'b0;
assign   tb_o_tag[18]                        =   tb_o_tag[17];

// CLK no. 19/1240
// *************************************************
assign   tb_i_valid[19]                      =   1'b0;
assign   tb_i_reset[19]                      =   1'b0;
assign   tb_i_sop[19]                        =   1'b0;
assign   tb_i_key_update[19]                 =   1'b0;
assign   tb_i_key[19]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[19]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[19]               =   1'b0;
assign   tb_i_rf_static_encrypt[19]          =   1'b1;
assign   tb_i_clear_fault_flags[19]          =   1'b0;
assign   tb_i_rf_static_aad_length[19]       =   64'h0000000000000100;
assign   tb_i_aad[19]                        =   tb_i_aad[18];
assign   tb_i_rf_static_plaintext_length[19] =   64'h0000000000000200;
assign   tb_i_plaintext[19]                  =   tb_i_plaintext[18];
assign   tb_o_valid[19]                      =   1'b0;
assign   tb_o_sop[19]                        =   1'b0;
assign   tb_o_ciphertext[19]                 =   tb_o_ciphertext[18];
assign   tb_o_tag_ready[19]                  =   1'b0;
assign   tb_o_tag[19]                        =   tb_o_tag[18];

// CLK no. 20/1240
// *************************************************
assign   tb_i_valid[20]                      =   1'b0;
assign   tb_i_reset[20]                      =   1'b0;
assign   tb_i_sop[20]                        =   1'b0;
assign   tb_i_key_update[20]                 =   1'b0;
assign   tb_i_key[20]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[20]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[20]               =   1'b0;
assign   tb_i_rf_static_encrypt[20]          =   1'b1;
assign   tb_i_clear_fault_flags[20]          =   1'b0;
assign   tb_i_rf_static_aad_length[20]       =   64'h0000000000000100;
assign   tb_i_aad[20]                        =   tb_i_aad[19];
assign   tb_i_rf_static_plaintext_length[20] =   64'h0000000000000200;
assign   tb_i_plaintext[20]                  =   tb_i_plaintext[19];
assign   tb_o_valid[20]                      =   1'b0;
assign   tb_o_sop[20]                        =   1'b0;
assign   tb_o_ciphertext[20]                 =   tb_o_ciphertext[19];
assign   tb_o_tag_ready[20]                  =   1'b0;
assign   tb_o_tag[20]                        =   tb_o_tag[19];

// CLK no. 21/1240
// *************************************************
assign   tb_i_valid[21]                      =   1'b0;
assign   tb_i_reset[21]                      =   1'b0;
assign   tb_i_sop[21]                        =   1'b0;
assign   tb_i_key_update[21]                 =   1'b0;
assign   tb_i_key[21]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[21]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[21]               =   1'b0;
assign   tb_i_rf_static_encrypt[21]          =   1'b1;
assign   tb_i_clear_fault_flags[21]          =   1'b0;
assign   tb_i_rf_static_aad_length[21]       =   64'h0000000000000100;
assign   tb_i_aad[21]                        =   tb_i_aad[20];
assign   tb_i_rf_static_plaintext_length[21] =   64'h0000000000000200;
assign   tb_i_plaintext[21]                  =   tb_i_plaintext[20];
assign   tb_o_valid[21]                      =   1'b0;
assign   tb_o_sop[21]                        =   1'b0;
assign   tb_o_ciphertext[21]                 =   tb_o_ciphertext[20];
assign   tb_o_tag_ready[21]                  =   1'b0;
assign   tb_o_tag[21]                        =   tb_o_tag[20];

// CLK no. 22/1240
// *************************************************
assign   tb_i_valid[22]                      =   1'b0;
assign   tb_i_reset[22]                      =   1'b0;
assign   tb_i_sop[22]                        =   1'b0;
assign   tb_i_key_update[22]                 =   1'b0;
assign   tb_i_key[22]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[22]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[22]               =   1'b0;
assign   tb_i_rf_static_encrypt[22]          =   1'b1;
assign   tb_i_clear_fault_flags[22]          =   1'b0;
assign   tb_i_rf_static_aad_length[22]       =   64'h0000000000000100;
assign   tb_i_aad[22]                        =   tb_i_aad[21];
assign   tb_i_rf_static_plaintext_length[22] =   64'h0000000000000200;
assign   tb_i_plaintext[22]                  =   tb_i_plaintext[21];
assign   tb_o_valid[22]                      =   1'b0;
assign   tb_o_sop[22]                        =   1'b0;
assign   tb_o_ciphertext[22]                 =   tb_o_ciphertext[21];
assign   tb_o_tag_ready[22]                  =   1'b0;
assign   tb_o_tag[22]                        =   tb_o_tag[21];

// CLK no. 23/1240
// *************************************************
assign   tb_i_valid[23]                      =   1'b0;
assign   tb_i_reset[23]                      =   1'b0;
assign   tb_i_sop[23]                        =   1'b0;
assign   tb_i_key_update[23]                 =   1'b0;
assign   tb_i_key[23]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[23]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[23]               =   1'b0;
assign   tb_i_rf_static_encrypt[23]          =   1'b1;
assign   tb_i_clear_fault_flags[23]          =   1'b0;
assign   tb_i_rf_static_aad_length[23]       =   64'h0000000000000100;
assign   tb_i_aad[23]                        =   tb_i_aad[22];
assign   tb_i_rf_static_plaintext_length[23] =   64'h0000000000000200;
assign   tb_i_plaintext[23]                  =   tb_i_plaintext[22];
assign   tb_o_valid[23]                      =   1'b0;
assign   tb_o_sop[23]                        =   1'b0;
assign   tb_o_ciphertext[23]                 =   tb_o_ciphertext[22];
assign   tb_o_tag_ready[23]                  =   1'b0;
assign   tb_o_tag[23]                        =   tb_o_tag[22];

// CLK no. 24/1240
// *************************************************
assign   tb_i_valid[24]                      =   1'b0;
assign   tb_i_reset[24]                      =   1'b0;
assign   tb_i_sop[24]                        =   1'b0;
assign   tb_i_key_update[24]                 =   1'b0;
assign   tb_i_key[24]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[24]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[24]               =   1'b0;
assign   tb_i_rf_static_encrypt[24]          =   1'b1;
assign   tb_i_clear_fault_flags[24]          =   1'b0;
assign   tb_i_rf_static_aad_length[24]       =   64'h0000000000000100;
assign   tb_i_aad[24]                        =   tb_i_aad[23];
assign   tb_i_rf_static_plaintext_length[24] =   64'h0000000000000200;
assign   tb_i_plaintext[24]                  =   tb_i_plaintext[23];
assign   tb_o_valid[24]                      =   1'b0;
assign   tb_o_sop[24]                        =   1'b0;
assign   tb_o_ciphertext[24]                 =   tb_o_ciphertext[23];
assign   tb_o_tag_ready[24]                  =   1'b0;
assign   tb_o_tag[24]                        =   tb_o_tag[23];

// CLK no. 25/1240
// *************************************************
assign   tb_i_valid[25]                      =   1'b0;
assign   tb_i_reset[25]                      =   1'b0;
assign   tb_i_sop[25]                        =   1'b0;
assign   tb_i_key_update[25]                 =   1'b0;
assign   tb_i_key[25]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[25]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[25]               =   1'b0;
assign   tb_i_rf_static_encrypt[25]          =   1'b1;
assign   tb_i_clear_fault_flags[25]          =   1'b0;
assign   tb_i_rf_static_aad_length[25]       =   64'h0000000000000100;
assign   tb_i_aad[25]                        =   tb_i_aad[24];
assign   tb_i_rf_static_plaintext_length[25] =   64'h0000000000000200;
assign   tb_i_plaintext[25]                  =   tb_i_plaintext[24];
assign   tb_o_valid[25]                      =   1'b0;
assign   tb_o_sop[25]                        =   1'b0;
assign   tb_o_ciphertext[25]                 =   tb_o_ciphertext[24];
assign   tb_o_tag_ready[25]                  =   1'b0;
assign   tb_o_tag[25]                        =   tb_o_tag[24];

// CLK no. 26/1240
// *************************************************
assign   tb_i_valid[26]                      =   1'b0;
assign   tb_i_reset[26]                      =   1'b0;
assign   tb_i_sop[26]                        =   1'b0;
assign   tb_i_key_update[26]                 =   1'b0;
assign   tb_i_key[26]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[26]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[26]               =   1'b0;
assign   tb_i_rf_static_encrypt[26]          =   1'b1;
assign   tb_i_clear_fault_flags[26]          =   1'b0;
assign   tb_i_rf_static_aad_length[26]       =   64'h0000000000000100;
assign   tb_i_aad[26]                        =   tb_i_aad[25];
assign   tb_i_rf_static_plaintext_length[26] =   64'h0000000000000200;
assign   tb_i_plaintext[26]                  =   tb_i_plaintext[25];
assign   tb_o_valid[26]                      =   1'b0;
assign   tb_o_sop[26]                        =   1'b0;
assign   tb_o_ciphertext[26]                 =   tb_o_ciphertext[25];
assign   tb_o_tag_ready[26]                  =   1'b0;
assign   tb_o_tag[26]                        =   tb_o_tag[25];

// CLK no. 27/1240
// *************************************************
assign   tb_i_valid[27]                      =   1'b0;
assign   tb_i_reset[27]                      =   1'b0;
assign   tb_i_sop[27]                        =   1'b0;
assign   tb_i_key_update[27]                 =   1'b0;
assign   tb_i_key[27]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[27]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[27]               =   1'b0;
assign   tb_i_rf_static_encrypt[27]          =   1'b1;
assign   tb_i_clear_fault_flags[27]          =   1'b0;
assign   tb_i_rf_static_aad_length[27]       =   64'h0000000000000100;
assign   tb_i_aad[27]                        =   tb_i_aad[26];
assign   tb_i_rf_static_plaintext_length[27] =   64'h0000000000000200;
assign   tb_i_plaintext[27]                  =   tb_i_plaintext[26];
assign   tb_o_valid[27]                      =   1'b0;
assign   tb_o_sop[27]                        =   1'b0;
assign   tb_o_ciphertext[27]                 =   tb_o_ciphertext[26];
assign   tb_o_tag_ready[27]                  =   1'b0;
assign   tb_o_tag[27]                        =   tb_o_tag[26];

// CLK no. 28/1240
// *************************************************
assign   tb_i_valid[28]                      =   1'b0;
assign   tb_i_reset[28]                      =   1'b0;
assign   tb_i_sop[28]                        =   1'b0;
assign   tb_i_key_update[28]                 =   1'b0;
assign   tb_i_key[28]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[28]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[28]               =   1'b0;
assign   tb_i_rf_static_encrypt[28]          =   1'b1;
assign   tb_i_clear_fault_flags[28]          =   1'b0;
assign   tb_i_rf_static_aad_length[28]       =   64'h0000000000000100;
assign   tb_i_aad[28]                        =   tb_i_aad[27];
assign   tb_i_rf_static_plaintext_length[28] =   64'h0000000000000200;
assign   tb_i_plaintext[28]                  =   tb_i_plaintext[27];
assign   tb_o_valid[28]                      =   1'b0;
assign   tb_o_sop[28]                        =   1'b0;
assign   tb_o_ciphertext[28]                 =   tb_o_ciphertext[27];
assign   tb_o_tag_ready[28]                  =   1'b0;
assign   tb_o_tag[28]                        =   tb_o_tag[27];

// CLK no. 29/1240
// *************************************************
assign   tb_i_valid[29]                      =   1'b0;
assign   tb_i_reset[29]                      =   1'b0;
assign   tb_i_sop[29]                        =   1'b0;
assign   tb_i_key_update[29]                 =   1'b0;
assign   tb_i_key[29]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[29]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[29]               =   1'b0;
assign   tb_i_rf_static_encrypt[29]          =   1'b1;
assign   tb_i_clear_fault_flags[29]          =   1'b0;
assign   tb_i_rf_static_aad_length[29]       =   64'h0000000000000100;
assign   tb_i_aad[29]                        =   tb_i_aad[28];
assign   tb_i_rf_static_plaintext_length[29] =   64'h0000000000000200;
assign   tb_i_plaintext[29]                  =   tb_i_plaintext[28];
assign   tb_o_valid[29]                      =   1'b0;
assign   tb_o_sop[29]                        =   1'b0;
assign   tb_o_ciphertext[29]                 =   tb_o_ciphertext[28];
assign   tb_o_tag_ready[29]                  =   1'b0;
assign   tb_o_tag[29]                        =   tb_o_tag[28];

// CLK no. 30/1240
// *************************************************
assign   tb_i_valid[30]                      =   1'b0;
assign   tb_i_reset[30]                      =   1'b0;
assign   tb_i_sop[30]                        =   1'b0;
assign   tb_i_key_update[30]                 =   1'b0;
assign   tb_i_key[30]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[30]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[30]               =   1'b0;
assign   tb_i_rf_static_encrypt[30]          =   1'b1;
assign   tb_i_clear_fault_flags[30]          =   1'b0;
assign   tb_i_rf_static_aad_length[30]       =   64'h0000000000000100;
assign   tb_i_aad[30]                        =   tb_i_aad[29];
assign   tb_i_rf_static_plaintext_length[30] =   64'h0000000000000200;
assign   tb_i_plaintext[30]                  =   tb_i_plaintext[29];
assign   tb_o_valid[30]                      =   1'b0;
assign   tb_o_sop[30]                        =   1'b0;
assign   tb_o_ciphertext[30]                 =   tb_o_ciphertext[29];
assign   tb_o_tag_ready[30]                  =   1'b0;
assign   tb_o_tag[30]                        =   tb_o_tag[29];

// CLK no. 31/1240
// *************************************************
assign   tb_i_valid[31]                      =   1'b0;
assign   tb_i_reset[31]                      =   1'b0;
assign   tb_i_sop[31]                        =   1'b0;
assign   tb_i_key_update[31]                 =   1'b0;
assign   tb_i_key[31]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[31]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[31]               =   1'b0;
assign   tb_i_rf_static_encrypt[31]          =   1'b1;
assign   tb_i_clear_fault_flags[31]          =   1'b0;
assign   tb_i_rf_static_aad_length[31]       =   64'h0000000000000100;
assign   tb_i_aad[31]                        =   tb_i_aad[30];
assign   tb_i_rf_static_plaintext_length[31] =   64'h0000000000000200;
assign   tb_i_plaintext[31]                  =   tb_i_plaintext[30];
assign   tb_o_valid[31]                      =   1'b0;
assign   tb_o_sop[31]                        =   1'b0;
assign   tb_o_ciphertext[31]                 =   tb_o_ciphertext[30];
assign   tb_o_tag_ready[31]                  =   1'b0;
assign   tb_o_tag[31]                        =   tb_o_tag[30];

// CLK no. 32/1240
// *************************************************
assign   tb_i_valid[32]                      =   1'b0;
assign   tb_i_reset[32]                      =   1'b0;
assign   tb_i_sop[32]                        =   1'b0;
assign   tb_i_key_update[32]                 =   1'b0;
assign   tb_i_key[32]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[32]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[32]               =   1'b0;
assign   tb_i_rf_static_encrypt[32]          =   1'b1;
assign   tb_i_clear_fault_flags[32]          =   1'b0;
assign   tb_i_rf_static_aad_length[32]       =   64'h0000000000000100;
assign   tb_i_aad[32]                        =   tb_i_aad[31];
assign   tb_i_rf_static_plaintext_length[32] =   64'h0000000000000200;
assign   tb_i_plaintext[32]                  =   tb_i_plaintext[31];
assign   tb_o_valid[32]                      =   1'b0;
assign   tb_o_sop[32]                        =   1'b0;
assign   tb_o_ciphertext[32]                 =   tb_o_ciphertext[31];
assign   tb_o_tag_ready[32]                  =   1'b0;
assign   tb_o_tag[32]                        =   tb_o_tag[31];

// CLK no. 33/1240
// *************************************************
assign   tb_i_valid[33]                      =   1'b0;
assign   tb_i_reset[33]                      =   1'b0;
assign   tb_i_sop[33]                        =   1'b0;
assign   tb_i_key_update[33]                 =   1'b0;
assign   tb_i_key[33]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[33]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[33]               =   1'b0;
assign   tb_i_rf_static_encrypt[33]          =   1'b1;
assign   tb_i_clear_fault_flags[33]          =   1'b0;
assign   tb_i_rf_static_aad_length[33]       =   64'h0000000000000100;
assign   tb_i_aad[33]                        =   tb_i_aad[32];
assign   tb_i_rf_static_plaintext_length[33] =   64'h0000000000000200;
assign   tb_i_plaintext[33]                  =   tb_i_plaintext[32];
assign   tb_o_valid[33]                      =   1'b0;
assign   tb_o_sop[33]                        =   1'b0;
assign   tb_o_ciphertext[33]                 =   tb_o_ciphertext[32];
assign   tb_o_tag_ready[33]                  =   1'b0;
assign   tb_o_tag[33]                        =   tb_o_tag[32];

// CLK no. 34/1240
// *************************************************
assign   tb_i_valid[34]                      =   1'b0;
assign   tb_i_reset[34]                      =   1'b0;
assign   tb_i_sop[34]                        =   1'b0;
assign   tb_i_key_update[34]                 =   1'b0;
assign   tb_i_key[34]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[34]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[34]               =   1'b0;
assign   tb_i_rf_static_encrypt[34]          =   1'b1;
assign   tb_i_clear_fault_flags[34]          =   1'b0;
assign   tb_i_rf_static_aad_length[34]       =   64'h0000000000000100;
assign   tb_i_aad[34]                        =   tb_i_aad[33];
assign   tb_i_rf_static_plaintext_length[34] =   64'h0000000000000200;
assign   tb_i_plaintext[34]                  =   tb_i_plaintext[33];
assign   tb_o_valid[34]                      =   1'b0;
assign   tb_o_sop[34]                        =   1'b0;
assign   tb_o_ciphertext[34]                 =   tb_o_ciphertext[33];
assign   tb_o_tag_ready[34]                  =   1'b0;
assign   tb_o_tag[34]                        =   tb_o_tag[33];

// CLK no. 35/1240
// *************************************************
assign   tb_i_valid[35]                      =   1'b0;
assign   tb_i_reset[35]                      =   1'b0;
assign   tb_i_sop[35]                        =   1'b0;
assign   tb_i_key_update[35]                 =   1'b0;
assign   tb_i_key[35]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[35]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[35]               =   1'b0;
assign   tb_i_rf_static_encrypt[35]          =   1'b1;
assign   tb_i_clear_fault_flags[35]          =   1'b0;
assign   tb_i_rf_static_aad_length[35]       =   64'h0000000000000100;
assign   tb_i_aad[35]                        =   tb_i_aad[34];
assign   tb_i_rf_static_plaintext_length[35] =   64'h0000000000000200;
assign   tb_i_plaintext[35]                  =   tb_i_plaintext[34];
assign   tb_o_valid[35]                      =   1'b0;
assign   tb_o_sop[35]                        =   1'b0;
assign   tb_o_ciphertext[35]                 =   tb_o_ciphertext[34];
assign   tb_o_tag_ready[35]                  =   1'b0;
assign   tb_o_tag[35]                        =   tb_o_tag[34];

// CLK no. 36/1240
// *************************************************
assign   tb_i_valid[36]                      =   1'b0;
assign   tb_i_reset[36]                      =   1'b0;
assign   tb_i_sop[36]                        =   1'b0;
assign   tb_i_key_update[36]                 =   1'b0;
assign   tb_i_key[36]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[36]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[36]               =   1'b0;
assign   tb_i_rf_static_encrypt[36]          =   1'b1;
assign   tb_i_clear_fault_flags[36]          =   1'b0;
assign   tb_i_rf_static_aad_length[36]       =   64'h0000000000000100;
assign   tb_i_aad[36]                        =   tb_i_aad[35];
assign   tb_i_rf_static_plaintext_length[36] =   64'h0000000000000200;
assign   tb_i_plaintext[36]                  =   tb_i_plaintext[35];
assign   tb_o_valid[36]                      =   1'b0;
assign   tb_o_sop[36]                        =   1'b0;
assign   tb_o_ciphertext[36]                 =   tb_o_ciphertext[35];
assign   tb_o_tag_ready[36]                  =   1'b0;
assign   tb_o_tag[36]                        =   tb_o_tag[35];

// CLK no. 37/1240
// *************************************************
assign   tb_i_valid[37]                      =   1'b0;
assign   tb_i_reset[37]                      =   1'b0;
assign   tb_i_sop[37]                        =   1'b0;
assign   tb_i_key_update[37]                 =   1'b0;
assign   tb_i_key[37]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[37]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[37]               =   1'b0;
assign   tb_i_rf_static_encrypt[37]          =   1'b1;
assign   tb_i_clear_fault_flags[37]          =   1'b0;
assign   tb_i_rf_static_aad_length[37]       =   64'h0000000000000100;
assign   tb_i_aad[37]                        =   tb_i_aad[36];
assign   tb_i_rf_static_plaintext_length[37] =   64'h0000000000000200;
assign   tb_i_plaintext[37]                  =   tb_i_plaintext[36];
assign   tb_o_valid[37]                      =   1'b0;
assign   tb_o_sop[37]                        =   1'b0;
assign   tb_o_ciphertext[37]                 =   tb_o_ciphertext[36];
assign   tb_o_tag_ready[37]                  =   1'b0;
assign   tb_o_tag[37]                        =   tb_o_tag[36];

// CLK no. 38/1240
// *************************************************
assign   tb_i_valid[38]                      =   1'b0;
assign   tb_i_reset[38]                      =   1'b0;
assign   tb_i_sop[38]                        =   1'b0;
assign   tb_i_key_update[38]                 =   1'b0;
assign   tb_i_key[38]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[38]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[38]               =   1'b0;
assign   tb_i_rf_static_encrypt[38]          =   1'b1;
assign   tb_i_clear_fault_flags[38]          =   1'b0;
assign   tb_i_rf_static_aad_length[38]       =   64'h0000000000000100;
assign   tb_i_aad[38]                        =   tb_i_aad[37];
assign   tb_i_rf_static_plaintext_length[38] =   64'h0000000000000200;
assign   tb_i_plaintext[38]                  =   tb_i_plaintext[37];
assign   tb_o_valid[38]                      =   1'b0;
assign   tb_o_sop[38]                        =   1'b0;
assign   tb_o_ciphertext[38]                 =   tb_o_ciphertext[37];
assign   tb_o_tag_ready[38]                  =   1'b0;
assign   tb_o_tag[38]                        =   tb_o_tag[37];

// CLK no. 39/1240
// *************************************************
assign   tb_i_valid[39]                      =   1'b0;
assign   tb_i_reset[39]                      =   1'b0;
assign   tb_i_sop[39]                        =   1'b0;
assign   tb_i_key_update[39]                 =   1'b0;
assign   tb_i_key[39]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[39]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[39]               =   1'b0;
assign   tb_i_rf_static_encrypt[39]          =   1'b1;
assign   tb_i_clear_fault_flags[39]          =   1'b0;
assign   tb_i_rf_static_aad_length[39]       =   64'h0000000000000100;
assign   tb_i_aad[39]                        =   tb_i_aad[38];
assign   tb_i_rf_static_plaintext_length[39] =   64'h0000000000000200;
assign   tb_i_plaintext[39]                  =   tb_i_plaintext[38];
assign   tb_o_valid[39]                      =   1'b0;
assign   tb_o_sop[39]                        =   1'b0;
assign   tb_o_ciphertext[39]                 =   tb_o_ciphertext[38];
assign   tb_o_tag_ready[39]                  =   1'b0;
assign   tb_o_tag[39]                        =   tb_o_tag[38];

// CLK no. 40/1240
// *************************************************
assign   tb_i_valid[40]                      =   1'b0;
assign   tb_i_reset[40]                      =   1'b0;
assign   tb_i_sop[40]                        =   1'b0;
assign   tb_i_key_update[40]                 =   1'b0;
assign   tb_i_key[40]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[40]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[40]               =   1'b0;
assign   tb_i_rf_static_encrypt[40]          =   1'b1;
assign   tb_i_clear_fault_flags[40]          =   1'b0;
assign   tb_i_rf_static_aad_length[40]       =   64'h0000000000000100;
assign   tb_i_aad[40]                        =   tb_i_aad[39];
assign   tb_i_rf_static_plaintext_length[40] =   64'h0000000000000200;
assign   tb_i_plaintext[40]                  =   tb_i_plaintext[39];
assign   tb_o_valid[40]                      =   1'b0;
assign   tb_o_sop[40]                        =   1'b0;
assign   tb_o_ciphertext[40]                 =   tb_o_ciphertext[39];
assign   tb_o_tag_ready[40]                  =   1'b0;
assign   tb_o_tag[40]                        =   tb_o_tag[39];

// CLK no. 41/1240
// *************************************************
assign   tb_i_valid[41]                      =   1'b0;
assign   tb_i_reset[41]                      =   1'b0;
assign   tb_i_sop[41]                        =   1'b0;
assign   tb_i_key_update[41]                 =   1'b0;
assign   tb_i_key[41]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[41]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[41]               =   1'b0;
assign   tb_i_rf_static_encrypt[41]          =   1'b1;
assign   tb_i_clear_fault_flags[41]          =   1'b0;
assign   tb_i_rf_static_aad_length[41]       =   64'h0000000000000100;
assign   tb_i_aad[41]                        =   tb_i_aad[40];
assign   tb_i_rf_static_plaintext_length[41] =   64'h0000000000000200;
assign   tb_i_plaintext[41]                  =   tb_i_plaintext[40];
assign   tb_o_valid[41]                      =   1'b0;
assign   tb_o_sop[41]                        =   1'b0;
assign   tb_o_ciphertext[41]                 =   tb_o_ciphertext[40];
assign   tb_o_tag_ready[41]                  =   1'b0;
assign   tb_o_tag[41]                        =   tb_o_tag[40];

// CLK no. 42/1240
// *************************************************
assign   tb_i_valid[42]                      =   1'b0;
assign   tb_i_reset[42]                      =   1'b0;
assign   tb_i_sop[42]                        =   1'b0;
assign   tb_i_key_update[42]                 =   1'b0;
assign   tb_i_key[42]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[42]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[42]               =   1'b0;
assign   tb_i_rf_static_encrypt[42]          =   1'b1;
assign   tb_i_clear_fault_flags[42]          =   1'b0;
assign   tb_i_rf_static_aad_length[42]       =   64'h0000000000000100;
assign   tb_i_aad[42]                        =   tb_i_aad[41];
assign   tb_i_rf_static_plaintext_length[42] =   64'h0000000000000200;
assign   tb_i_plaintext[42]                  =   tb_i_plaintext[41];
assign   tb_o_valid[42]                      =   1'b0;
assign   tb_o_sop[42]                        =   1'b0;
assign   tb_o_ciphertext[42]                 =   tb_o_ciphertext[41];
assign   tb_o_tag_ready[42]                  =   1'b0;
assign   tb_o_tag[42]                        =   tb_o_tag[41];

// CLK no. 43/1240
// *************************************************
assign   tb_i_valid[43]                      =   1'b0;
assign   tb_i_reset[43]                      =   1'b0;
assign   tb_i_sop[43]                        =   1'b0;
assign   tb_i_key_update[43]                 =   1'b0;
assign   tb_i_key[43]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[43]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[43]               =   1'b0;
assign   tb_i_rf_static_encrypt[43]          =   1'b1;
assign   tb_i_clear_fault_flags[43]          =   1'b0;
assign   tb_i_rf_static_aad_length[43]       =   64'h0000000000000100;
assign   tb_i_aad[43]                        =   tb_i_aad[42];
assign   tb_i_rf_static_plaintext_length[43] =   64'h0000000000000200;
assign   tb_i_plaintext[43]                  =   tb_i_plaintext[42];
assign   tb_o_valid[43]                      =   1'b0;
assign   tb_o_sop[43]                        =   1'b0;
assign   tb_o_ciphertext[43]                 =   tb_o_ciphertext[42];
assign   tb_o_tag_ready[43]                  =   1'b0;
assign   tb_o_tag[43]                        =   tb_o_tag[42];

// CLK no. 44/1240
// *************************************************
assign   tb_i_valid[44]                      =   1'b0;
assign   tb_i_reset[44]                      =   1'b0;
assign   tb_i_sop[44]                        =   1'b0;
assign   tb_i_key_update[44]                 =   1'b0;
assign   tb_i_key[44]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[44]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[44]               =   1'b0;
assign   tb_i_rf_static_encrypt[44]          =   1'b1;
assign   tb_i_clear_fault_flags[44]          =   1'b0;
assign   tb_i_rf_static_aad_length[44]       =   64'h0000000000000100;
assign   tb_i_aad[44]                        =   tb_i_aad[43];
assign   tb_i_rf_static_plaintext_length[44] =   64'h0000000000000200;
assign   tb_i_plaintext[44]                  =   tb_i_plaintext[43];
assign   tb_o_valid[44]                      =   1'b0;
assign   tb_o_sop[44]                        =   1'b0;
assign   tb_o_ciphertext[44]                 =   tb_o_ciphertext[43];
assign   tb_o_tag_ready[44]                  =   1'b0;
assign   tb_o_tag[44]                        =   tb_o_tag[43];

// CLK no. 45/1240
// *************************************************
assign   tb_i_valid[45]                      =   1'b0;
assign   tb_i_reset[45]                      =   1'b0;
assign   tb_i_sop[45]                        =   1'b0;
assign   tb_i_key_update[45]                 =   1'b0;
assign   tb_i_key[45]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[45]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[45]               =   1'b0;
assign   tb_i_rf_static_encrypt[45]          =   1'b1;
assign   tb_i_clear_fault_flags[45]          =   1'b0;
assign   tb_i_rf_static_aad_length[45]       =   64'h0000000000000100;
assign   tb_i_aad[45]                        =   tb_i_aad[44];
assign   tb_i_rf_static_plaintext_length[45] =   64'h0000000000000200;
assign   tb_i_plaintext[45]                  =   tb_i_plaintext[44];
assign   tb_o_valid[45]                      =   1'b0;
assign   tb_o_sop[45]                        =   1'b0;
assign   tb_o_ciphertext[45]                 =   tb_o_ciphertext[44];
assign   tb_o_tag_ready[45]                  =   1'b0;
assign   tb_o_tag[45]                        =   tb_o_tag[44];

// CLK no. 46/1240
// *************************************************
assign   tb_i_valid[46]                      =   1'b0;
assign   tb_i_reset[46]                      =   1'b0;
assign   tb_i_sop[46]                        =   1'b0;
assign   tb_i_key_update[46]                 =   1'b0;
assign   tb_i_key[46]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[46]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[46]               =   1'b0;
assign   tb_i_rf_static_encrypt[46]          =   1'b1;
assign   tb_i_clear_fault_flags[46]          =   1'b0;
assign   tb_i_rf_static_aad_length[46]       =   64'h0000000000000100;
assign   tb_i_aad[46]                        =   tb_i_aad[45];
assign   tb_i_rf_static_plaintext_length[46] =   64'h0000000000000200;
assign   tb_i_plaintext[46]                  =   tb_i_plaintext[45];
assign   tb_o_valid[46]                      =   1'b0;
assign   tb_o_sop[46]                        =   1'b0;
assign   tb_o_ciphertext[46]                 =   tb_o_ciphertext[45];
assign   tb_o_tag_ready[46]                  =   1'b0;
assign   tb_o_tag[46]                        =   tb_o_tag[45];

// CLK no. 47/1240
// *************************************************
assign   tb_i_valid[47]                      =   1'b0;
assign   tb_i_reset[47]                      =   1'b0;
assign   tb_i_sop[47]                        =   1'b0;
assign   tb_i_key_update[47]                 =   1'b0;
assign   tb_i_key[47]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[47]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[47]               =   1'b0;
assign   tb_i_rf_static_encrypt[47]          =   1'b1;
assign   tb_i_clear_fault_flags[47]          =   1'b0;
assign   tb_i_rf_static_aad_length[47]       =   64'h0000000000000100;
assign   tb_i_aad[47]                        =   tb_i_aad[46];
assign   tb_i_rf_static_plaintext_length[47] =   64'h0000000000000200;
assign   tb_i_plaintext[47]                  =   tb_i_plaintext[46];
assign   tb_o_valid[47]                      =   1'b1;
assign   tb_o_sop[47]                        =   1'b1;
assign   tb_o_ciphertext[47]                 =   256'h5d1ea585cded914114b5d5f8b1abde5288c1e0dc6fa60d49200577b4406e873b;
assign   tb_o_tag_ready[47]                  =   1'b0;
assign   tb_o_tag[47]                        =   tb_o_tag[46];

// CLK no. 48/1240
// *************************************************
assign   tb_i_valid[48]                      =   1'b0;
assign   tb_i_reset[48]                      =   1'b0;
assign   tb_i_sop[48]                        =   1'b0;
assign   tb_i_key_update[48]                 =   1'b0;
assign   tb_i_key[48]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[48]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[48]               =   1'b0;
assign   tb_i_rf_static_encrypt[48]          =   1'b1;
assign   tb_i_clear_fault_flags[48]          =   1'b0;
assign   tb_i_rf_static_aad_length[48]       =   64'h0000000000000100;
assign   tb_i_aad[48]                        =   tb_i_aad[47];
assign   tb_i_rf_static_plaintext_length[48] =   64'h0000000000000200;
assign   tb_i_plaintext[48]                  =   tb_i_plaintext[47];
assign   tb_o_valid[48]                      =   1'b1;
assign   tb_o_sop[48]                        =   1'b0;
assign   tb_o_ciphertext[48]                 =   256'h7df9caf3ff7c8c744d242bbb07a088c46fc0a9bf5f74178ec7a3174d0e3bf095;
assign   tb_o_tag_ready[48]                  =   1'b0;
assign   tb_o_tag[48]                        =   tb_o_tag[47];

// CLK no. 49/1240
// *************************************************
assign   tb_i_valid[49]                      =   1'b0;
assign   tb_i_reset[49]                      =   1'b0;
assign   tb_i_sop[49]                        =   1'b0;
assign   tb_i_key_update[49]                 =   1'b0;
assign   tb_i_key[49]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[49]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[49]               =   1'b0;
assign   tb_i_rf_static_encrypt[49]          =   1'b1;
assign   tb_i_clear_fault_flags[49]          =   1'b0;
assign   tb_i_rf_static_aad_length[49]       =   64'h0000000000000100;
assign   tb_i_aad[49]                        =   tb_i_aad[48];
assign   tb_i_rf_static_plaintext_length[49] =   64'h0000000000000200;
assign   tb_i_plaintext[49]                  =   tb_i_plaintext[48];
assign   tb_o_valid[49]                      =   1'b0;
assign   tb_o_sop[49]                        =   1'b0;
assign   tb_o_ciphertext[49]                 =   tb_o_ciphertext[48];
assign   tb_o_tag_ready[49]                  =   1'b0;
assign   tb_o_tag[49]                        =   tb_o_tag[48];

// CLK no. 50/1240
// *************************************************
assign   tb_i_valid[50]                      =   1'b0;
assign   tb_i_reset[50]                      =   1'b0;
assign   tb_i_sop[50]                        =   1'b0;
assign   tb_i_key_update[50]                 =   1'b0;
assign   tb_i_key[50]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[50]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[50]               =   1'b0;
assign   tb_i_rf_static_encrypt[50]          =   1'b1;
assign   tb_i_clear_fault_flags[50]          =   1'b0;
assign   tb_i_rf_static_aad_length[50]       =   64'h0000000000000100;
assign   tb_i_aad[50]                        =   tb_i_aad[49];
assign   tb_i_rf_static_plaintext_length[50] =   64'h0000000000000200;
assign   tb_i_plaintext[50]                  =   tb_i_plaintext[49];
assign   tb_o_valid[50]                      =   1'b0;
assign   tb_o_sop[50]                        =   1'b0;
assign   tb_o_ciphertext[50]                 =   tb_o_ciphertext[49];
assign   tb_o_tag_ready[50]                  =   1'b0;
assign   tb_o_tag[50]                        =   tb_o_tag[49];

// CLK no. 51/1240
// *************************************************
assign   tb_i_valid[51]                      =   1'b0;
assign   tb_i_reset[51]                      =   1'b0;
assign   tb_i_sop[51]                        =   1'b0;
assign   tb_i_key_update[51]                 =   1'b0;
assign   tb_i_key[51]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[51]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[51]               =   1'b0;
assign   tb_i_rf_static_encrypt[51]          =   1'b1;
assign   tb_i_clear_fault_flags[51]          =   1'b0;
assign   tb_i_rf_static_aad_length[51]       =   64'h0000000000000100;
assign   tb_i_aad[51]                        =   tb_i_aad[50];
assign   tb_i_rf_static_plaintext_length[51] =   64'h0000000000000200;
assign   tb_i_plaintext[51]                  =   tb_i_plaintext[50];
assign   tb_o_valid[51]                      =   1'b0;
assign   tb_o_sop[51]                        =   1'b0;
assign   tb_o_ciphertext[51]                 =   tb_o_ciphertext[50];
assign   tb_o_tag_ready[51]                  =   1'b0;
assign   tb_o_tag[51]                        =   tb_o_tag[50];

// CLK no. 52/1240
// *************************************************
assign   tb_i_valid[52]                      =   1'b0;
assign   tb_i_reset[52]                      =   1'b0;
assign   tb_i_sop[52]                        =   1'b0;
assign   tb_i_key_update[52]                 =   1'b0;
assign   tb_i_key[52]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[52]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[52]               =   1'b0;
assign   tb_i_rf_static_encrypt[52]          =   1'b1;
assign   tb_i_clear_fault_flags[52]          =   1'b0;
assign   tb_i_rf_static_aad_length[52]       =   64'h0000000000000100;
assign   tb_i_aad[52]                        =   tb_i_aad[51];
assign   tb_i_rf_static_plaintext_length[52] =   64'h0000000000000200;
assign   tb_i_plaintext[52]                  =   tb_i_plaintext[51];
assign   tb_o_valid[52]                      =   1'b0;
assign   tb_o_sop[52]                        =   1'b0;
assign   tb_o_ciphertext[52]                 =   tb_o_ciphertext[51];
assign   tb_o_tag_ready[52]                  =   1'b0;
assign   tb_o_tag[52]                        =   tb_o_tag[51];

// CLK no. 53/1240
// *************************************************
assign   tb_i_valid[53]                      =   1'b0;
assign   tb_i_reset[53]                      =   1'b0;
assign   tb_i_sop[53]                        =   1'b0;
assign   tb_i_key_update[53]                 =   1'b0;
assign   tb_i_key[53]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[53]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[53]               =   1'b0;
assign   tb_i_rf_static_encrypt[53]          =   1'b1;
assign   tb_i_clear_fault_flags[53]          =   1'b0;
assign   tb_i_rf_static_aad_length[53]       =   64'h0000000000000100;
assign   tb_i_aad[53]                        =   tb_i_aad[52];
assign   tb_i_rf_static_plaintext_length[53] =   64'h0000000000000200;
assign   tb_i_plaintext[53]                  =   tb_i_plaintext[52];
assign   tb_o_valid[53]                      =   1'b0;
assign   tb_o_sop[53]                        =   1'b0;
assign   tb_o_ciphertext[53]                 =   tb_o_ciphertext[52];
assign   tb_o_tag_ready[53]                  =   1'b0;
assign   tb_o_tag[53]                        =   tb_o_tag[52];

// CLK no. 54/1240
// *************************************************
assign   tb_i_valid[54]                      =   1'b0;
assign   tb_i_reset[54]                      =   1'b0;
assign   tb_i_sop[54]                        =   1'b0;
assign   tb_i_key_update[54]                 =   1'b0;
assign   tb_i_key[54]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[54]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[54]               =   1'b0;
assign   tb_i_rf_static_encrypt[54]          =   1'b1;
assign   tb_i_clear_fault_flags[54]          =   1'b0;
assign   tb_i_rf_static_aad_length[54]       =   64'h0000000000000100;
assign   tb_i_aad[54]                        =   tb_i_aad[53];
assign   tb_i_rf_static_plaintext_length[54] =   64'h0000000000000200;
assign   tb_i_plaintext[54]                  =   tb_i_plaintext[53];
assign   tb_o_valid[54]                      =   1'b0;
assign   tb_o_sop[54]                        =   1'b0;
assign   tb_o_ciphertext[54]                 =   tb_o_ciphertext[53];
assign   tb_o_tag_ready[54]                  =   1'b0;
assign   tb_o_tag[54]                        =   tb_o_tag[53];

// CLK no. 55/1240
// *************************************************
assign   tb_i_valid[55]                      =   1'b0;
assign   tb_i_reset[55]                      =   1'b0;
assign   tb_i_sop[55]                        =   1'b0;
assign   tb_i_key_update[55]                 =   1'b0;
assign   tb_i_key[55]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[55]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[55]               =   1'b0;
assign   tb_i_rf_static_encrypt[55]          =   1'b1;
assign   tb_i_clear_fault_flags[55]          =   1'b0;
assign   tb_i_rf_static_aad_length[55]       =   64'h0000000000000100;
assign   tb_i_aad[55]                        =   tb_i_aad[54];
assign   tb_i_rf_static_plaintext_length[55] =   64'h0000000000000200;
assign   tb_i_plaintext[55]                  =   tb_i_plaintext[54];
assign   tb_o_valid[55]                      =   1'b0;
assign   tb_o_sop[55]                        =   1'b0;
assign   tb_o_ciphertext[55]                 =   tb_o_ciphertext[54];
assign   tb_o_tag_ready[55]                  =   1'b0;
assign   tb_o_tag[55]                        =   tb_o_tag[54];

// CLK no. 56/1240
// *************************************************
assign   tb_i_valid[56]                      =   1'b0;
assign   tb_i_reset[56]                      =   1'b0;
assign   tb_i_sop[56]                        =   1'b0;
assign   tb_i_key_update[56]                 =   1'b0;
assign   tb_i_key[56]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[56]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[56]               =   1'b0;
assign   tb_i_rf_static_encrypt[56]          =   1'b1;
assign   tb_i_clear_fault_flags[56]          =   1'b0;
assign   tb_i_rf_static_aad_length[56]       =   64'h0000000000000100;
assign   tb_i_aad[56]                        =   tb_i_aad[55];
assign   tb_i_rf_static_plaintext_length[56] =   64'h0000000000000200;
assign   tb_i_plaintext[56]                  =   tb_i_plaintext[55];
assign   tb_o_valid[56]                      =   1'b0;
assign   tb_o_sop[56]                        =   1'b0;
assign   tb_o_ciphertext[56]                 =   tb_o_ciphertext[55];
assign   tb_o_tag_ready[56]                  =   1'b0;
assign   tb_o_tag[56]                        =   tb_o_tag[55];

// CLK no. 57/1240
// *************************************************
assign   tb_i_valid[57]                      =   1'b0;
assign   tb_i_reset[57]                      =   1'b0;
assign   tb_i_sop[57]                        =   1'b0;
assign   tb_i_key_update[57]                 =   1'b0;
assign   tb_i_key[57]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[57]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[57]               =   1'b0;
assign   tb_i_rf_static_encrypt[57]          =   1'b1;
assign   tb_i_clear_fault_flags[57]          =   1'b0;
assign   tb_i_rf_static_aad_length[57]       =   64'h0000000000000100;
assign   tb_i_aad[57]                        =   tb_i_aad[56];
assign   tb_i_rf_static_plaintext_length[57] =   64'h0000000000000200;
assign   tb_i_plaintext[57]                  =   tb_i_plaintext[56];
assign   tb_o_valid[57]                      =   1'b0;
assign   tb_o_sop[57]                        =   1'b0;
assign   tb_o_ciphertext[57]                 =   tb_o_ciphertext[56];
assign   tb_o_tag_ready[57]                  =   1'b1;
assign   tb_o_tag[57]                        =   128'h5a915104103e269ed22e1f0beea00a8f;

// CLK no. 58/1240
// *************************************************
assign   tb_i_valid[58]                      =   1'b0;
assign   tb_i_reset[58]                      =   1'b0;
assign   tb_i_sop[58]                        =   1'b0;
assign   tb_i_key_update[58]                 =   1'b0;
assign   tb_i_key[58]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[58]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[58]               =   1'b0;
assign   tb_i_rf_static_encrypt[58]          =   1'b1;
assign   tb_i_clear_fault_flags[58]          =   1'b0;
assign   tb_i_rf_static_aad_length[58]       =   64'h0000000000000100;
assign   tb_i_aad[58]                        =   tb_i_aad[57];
assign   tb_i_rf_static_plaintext_length[58] =   64'h0000000000000200;
assign   tb_i_plaintext[58]                  =   tb_i_plaintext[57];
assign   tb_o_valid[58]                      =   1'b0;
assign   tb_o_sop[58]                        =   1'b0;
assign   tb_o_ciphertext[58]                 =   tb_o_ciphertext[57];
assign   tb_o_tag_ready[58]                  =   1'b0;
assign   tb_o_tag[58]                        =   tb_o_tag[57];

// CLK no. 59/1240
// *************************************************
assign   tb_i_valid[59]                      =   1'b0;
assign   tb_i_reset[59]                      =   1'b0;
assign   tb_i_sop[59]                        =   1'b0;
assign   tb_i_key_update[59]                 =   1'b0;
assign   tb_i_key[59]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[59]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[59]               =   1'b0;
assign   tb_i_rf_static_encrypt[59]          =   1'b1;
assign   tb_i_clear_fault_flags[59]          =   1'b0;
assign   tb_i_rf_static_aad_length[59]       =   64'h0000000000000100;
assign   tb_i_aad[59]                        =   tb_i_aad[58];
assign   tb_i_rf_static_plaintext_length[59] =   64'h0000000000000200;
assign   tb_i_plaintext[59]                  =   tb_i_plaintext[58];
assign   tb_o_valid[59]                      =   1'b0;
assign   tb_o_sop[59]                        =   1'b0;
assign   tb_o_ciphertext[59]                 =   tb_o_ciphertext[58];
assign   tb_o_tag_ready[59]                  =   1'b0;
assign   tb_o_tag[59]                        =   tb_o_tag[58];

// CLK no. 60/1240
// *************************************************
assign   tb_i_valid[60]                      =   1'b0;
assign   tb_i_reset[60]                      =   1'b0;
assign   tb_i_sop[60]                        =   1'b1;
assign   tb_i_key_update[60]                 =   1'b0;
assign   tb_i_key[60]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[60]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[60]               =   1'b0;
assign   tb_i_rf_static_encrypt[60]          =   1'b1;
assign   tb_i_clear_fault_flags[60]          =   1'b0;
assign   tb_i_rf_static_aad_length[60]       =   64'h0000000000000100;
assign   tb_i_aad[60]                        =   tb_i_aad[59];
assign   tb_i_rf_static_plaintext_length[60] =   64'h0000000000000280;
assign   tb_i_plaintext[60]                  =   tb_i_plaintext[59];
assign   tb_o_valid[60]                      =   1'b0;
assign   tb_o_sop[60]                        =   1'b0;
assign   tb_o_ciphertext[60]                 =   tb_o_ciphertext[59];
assign   tb_o_tag_ready[60]                  =   1'b0;
assign   tb_o_tag[60]                        =   tb_o_tag[59];

// CLK no. 61/1240
// *************************************************
assign   tb_i_valid[61]                      =   1'b1;
assign   tb_i_reset[61]                      =   1'b0;
assign   tb_i_sop[61]                        =   1'b0;
assign   tb_i_key_update[61]                 =   1'b0;
assign   tb_i_key[61]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[61]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[61]               =   1'b0;
assign   tb_i_rf_static_encrypt[61]          =   1'b1;
assign   tb_i_clear_fault_flags[61]          =   1'b0;
assign   tb_i_rf_static_aad_length[61]       =   64'h0000000000000100;
assign   tb_i_aad[61]                        =   256'h4229ca6bea2f24a558ab32d80601d879c3a378f03309a9c20a919c263b586311;
assign   tb_i_rf_static_plaintext_length[61] =   64'h0000000000000280;
assign   tb_i_plaintext[61]                  =   tb_i_plaintext[60];
assign   tb_o_valid[61]                      =   1'b0;
assign   tb_o_sop[61]                        =   1'b0;
assign   tb_o_ciphertext[61]                 =   tb_o_ciphertext[60];
assign   tb_o_tag_ready[61]                  =   1'b0;
assign   tb_o_tag[61]                        =   tb_o_tag[60];

// CLK no. 62/1240
// *************************************************
assign   tb_i_valid[62]                      =   1'b1;
assign   tb_i_reset[62]                      =   1'b0;
assign   tb_i_sop[62]                        =   1'b0;
assign   tb_i_key_update[62]                 =   1'b0;
assign   tb_i_key[62]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[62]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[62]               =   1'b0;
assign   tb_i_rf_static_encrypt[62]          =   1'b1;
assign   tb_i_clear_fault_flags[62]          =   1'b0;
assign   tb_i_rf_static_aad_length[62]       =   64'h0000000000000100;
assign   tb_i_aad[62]                        =   tb_i_aad[61];
assign   tb_i_rf_static_plaintext_length[62] =   64'h0000000000000280;
assign   tb_i_plaintext[62]                  =   256'hdfaa5d32397bcf2ef7577af6d3a067029be36fa8de79b621b6fea204e02e1f51;
assign   tb_o_valid[62]                      =   1'b0;
assign   tb_o_sop[62]                        =   1'b0;
assign   tb_o_ciphertext[62]                 =   tb_o_ciphertext[61];
assign   tb_o_tag_ready[62]                  =   1'b0;
assign   tb_o_tag[62]                        =   tb_o_tag[61];

// CLK no. 63/1240
// *************************************************
assign   tb_i_valid[63]                      =   1'b1;
assign   tb_i_reset[63]                      =   1'b0;
assign   tb_i_sop[63]                        =   1'b0;
assign   tb_i_key_update[63]                 =   1'b0;
assign   tb_i_key[63]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[63]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[63]               =   1'b0;
assign   tb_i_rf_static_encrypt[63]          =   1'b1;
assign   tb_i_clear_fault_flags[63]          =   1'b0;
assign   tb_i_rf_static_aad_length[63]       =   64'h0000000000000100;
assign   tb_i_aad[63]                        =   tb_i_aad[62];
assign   tb_i_rf_static_plaintext_length[63] =   64'h0000000000000280;
assign   tb_i_plaintext[63]                  =   256'hdf79ae285b5e9c052e66a68df6de90ffe378cacba44d3b8f17335f3304766e23;
assign   tb_o_valid[63]                      =   1'b0;
assign   tb_o_sop[63]                        =   1'b0;
assign   tb_o_ciphertext[63]                 =   tb_o_ciphertext[62];
assign   tb_o_tag_ready[63]                  =   1'b0;
assign   tb_o_tag[63]                        =   tb_o_tag[62];

// CLK no. 64/1240
// *************************************************
assign   tb_i_valid[64]                      =   1'b1;
assign   tb_i_reset[64]                      =   1'b0;
assign   tb_i_sop[64]                        =   1'b0;
assign   tb_i_key_update[64]                 =   1'b0;
assign   tb_i_key[64]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[64]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[64]               =   1'b0;
assign   tb_i_rf_static_encrypt[64]          =   1'b1;
assign   tb_i_clear_fault_flags[64]          =   1'b0;
assign   tb_i_rf_static_aad_length[64]       =   64'h0000000000000100;
assign   tb_i_aad[64]                        =   tb_i_aad[63];
assign   tb_i_rf_static_plaintext_length[64] =   64'h0000000000000280;
assign   tb_i_plaintext[64]                  =   256'h788b4279cf5f9af78ff906ca1f312d7b;
assign   tb_o_valid[64]                      =   1'b0;
assign   tb_o_sop[64]                        =   1'b0;
assign   tb_o_ciphertext[64]                 =   tb_o_ciphertext[63];
assign   tb_o_tag_ready[64]                  =   1'b0;
assign   tb_o_tag[64]                        =   tb_o_tag[63];

// CLK no. 65/1240
// *************************************************
assign   tb_i_valid[65]                      =   1'b0;
assign   tb_i_reset[65]                      =   1'b0;
assign   tb_i_sop[65]                        =   1'b0;
assign   tb_i_key_update[65]                 =   1'b0;
assign   tb_i_key[65]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[65]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[65]               =   1'b0;
assign   tb_i_rf_static_encrypt[65]          =   1'b1;
assign   tb_i_clear_fault_flags[65]          =   1'b0;
assign   tb_i_rf_static_aad_length[65]       =   64'h0000000000000100;
assign   tb_i_aad[65]                        =   tb_i_aad[64];
assign   tb_i_rf_static_plaintext_length[65] =   64'h0000000000000280;
assign   tb_i_plaintext[65]                  =   tb_i_plaintext[64];
assign   tb_o_valid[65]                      =   1'b0;
assign   tb_o_sop[65]                        =   1'b0;
assign   tb_o_ciphertext[65]                 =   tb_o_ciphertext[64];
assign   tb_o_tag_ready[65]                  =   1'b0;
assign   tb_o_tag[65]                        =   tb_o_tag[64];

// CLK no. 66/1240
// *************************************************
assign   tb_i_valid[66]                      =   1'b0;
assign   tb_i_reset[66]                      =   1'b0;
assign   tb_i_sop[66]                        =   1'b0;
assign   tb_i_key_update[66]                 =   1'b0;
assign   tb_i_key[66]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[66]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[66]               =   1'b0;
assign   tb_i_rf_static_encrypt[66]          =   1'b1;
assign   tb_i_clear_fault_flags[66]          =   1'b0;
assign   tb_i_rf_static_aad_length[66]       =   64'h0000000000000100;
assign   tb_i_aad[66]                        =   tb_i_aad[65];
assign   tb_i_rf_static_plaintext_length[66] =   64'h0000000000000280;
assign   tb_i_plaintext[66]                  =   tb_i_plaintext[65];
assign   tb_o_valid[66]                      =   1'b0;
assign   tb_o_sop[66]                        =   1'b0;
assign   tb_o_ciphertext[66]                 =   tb_o_ciphertext[65];
assign   tb_o_tag_ready[66]                  =   1'b0;
assign   tb_o_tag[66]                        =   tb_o_tag[65];

// CLK no. 67/1240
// *************************************************
assign   tb_i_valid[67]                      =   1'b0;
assign   tb_i_reset[67]                      =   1'b0;
assign   tb_i_sop[67]                        =   1'b0;
assign   tb_i_key_update[67]                 =   1'b0;
assign   tb_i_key[67]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[67]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[67]               =   1'b0;
assign   tb_i_rf_static_encrypt[67]          =   1'b1;
assign   tb_i_clear_fault_flags[67]          =   1'b0;
assign   tb_i_rf_static_aad_length[67]       =   64'h0000000000000100;
assign   tb_i_aad[67]                        =   tb_i_aad[66];
assign   tb_i_rf_static_plaintext_length[67] =   64'h0000000000000280;
assign   tb_i_plaintext[67]                  =   tb_i_plaintext[66];
assign   tb_o_valid[67]                      =   1'b0;
assign   tb_o_sop[67]                        =   1'b0;
assign   tb_o_ciphertext[67]                 =   tb_o_ciphertext[66];
assign   tb_o_tag_ready[67]                  =   1'b0;
assign   tb_o_tag[67]                        =   tb_o_tag[66];

// CLK no. 68/1240
// *************************************************
assign   tb_i_valid[68]                      =   1'b0;
assign   tb_i_reset[68]                      =   1'b0;
assign   tb_i_sop[68]                        =   1'b0;
assign   tb_i_key_update[68]                 =   1'b0;
assign   tb_i_key[68]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[68]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[68]               =   1'b0;
assign   tb_i_rf_static_encrypt[68]          =   1'b1;
assign   tb_i_clear_fault_flags[68]          =   1'b0;
assign   tb_i_rf_static_aad_length[68]       =   64'h0000000000000100;
assign   tb_i_aad[68]                        =   tb_i_aad[67];
assign   tb_i_rf_static_plaintext_length[68] =   64'h0000000000000280;
assign   tb_i_plaintext[68]                  =   tb_i_plaintext[67];
assign   tb_o_valid[68]                      =   1'b0;
assign   tb_o_sop[68]                        =   1'b0;
assign   tb_o_ciphertext[68]                 =   tb_o_ciphertext[67];
assign   tb_o_tag_ready[68]                  =   1'b0;
assign   tb_o_tag[68]                        =   tb_o_tag[67];

// CLK no. 69/1240
// *************************************************
assign   tb_i_valid[69]                      =   1'b0;
assign   tb_i_reset[69]                      =   1'b0;
assign   tb_i_sop[69]                        =   1'b0;
assign   tb_i_key_update[69]                 =   1'b0;
assign   tb_i_key[69]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[69]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[69]               =   1'b0;
assign   tb_i_rf_static_encrypt[69]          =   1'b1;
assign   tb_i_clear_fault_flags[69]          =   1'b0;
assign   tb_i_rf_static_aad_length[69]       =   64'h0000000000000100;
assign   tb_i_aad[69]                        =   tb_i_aad[68];
assign   tb_i_rf_static_plaintext_length[69] =   64'h0000000000000280;
assign   tb_i_plaintext[69]                  =   tb_i_plaintext[68];
assign   tb_o_valid[69]                      =   1'b0;
assign   tb_o_sop[69]                        =   1'b0;
assign   tb_o_ciphertext[69]                 =   tb_o_ciphertext[68];
assign   tb_o_tag_ready[69]                  =   1'b0;
assign   tb_o_tag[69]                        =   tb_o_tag[68];

// CLK no. 70/1240
// *************************************************
assign   tb_i_valid[70]                      =   1'b0;
assign   tb_i_reset[70]                      =   1'b0;
assign   tb_i_sop[70]                        =   1'b0;
assign   tb_i_key_update[70]                 =   1'b0;
assign   tb_i_key[70]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[70]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[70]               =   1'b0;
assign   tb_i_rf_static_encrypt[70]          =   1'b1;
assign   tb_i_clear_fault_flags[70]          =   1'b0;
assign   tb_i_rf_static_aad_length[70]       =   64'h0000000000000100;
assign   tb_i_aad[70]                        =   tb_i_aad[69];
assign   tb_i_rf_static_plaintext_length[70] =   64'h0000000000000280;
assign   tb_i_plaintext[70]                  =   tb_i_plaintext[69];
assign   tb_o_valid[70]                      =   1'b0;
assign   tb_o_sop[70]                        =   1'b0;
assign   tb_o_ciphertext[70]                 =   tb_o_ciphertext[69];
assign   tb_o_tag_ready[70]                  =   1'b0;
assign   tb_o_tag[70]                        =   tb_o_tag[69];

// CLK no. 71/1240
// *************************************************
assign   tb_i_valid[71]                      =   1'b0;
assign   tb_i_reset[71]                      =   1'b0;
assign   tb_i_sop[71]                        =   1'b0;
assign   tb_i_key_update[71]                 =   1'b0;
assign   tb_i_key[71]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[71]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[71]               =   1'b0;
assign   tb_i_rf_static_encrypt[71]          =   1'b1;
assign   tb_i_clear_fault_flags[71]          =   1'b0;
assign   tb_i_rf_static_aad_length[71]       =   64'h0000000000000100;
assign   tb_i_aad[71]                        =   tb_i_aad[70];
assign   tb_i_rf_static_plaintext_length[71] =   64'h0000000000000280;
assign   tb_i_plaintext[71]                  =   tb_i_plaintext[70];
assign   tb_o_valid[71]                      =   1'b0;
assign   tb_o_sop[71]                        =   1'b0;
assign   tb_o_ciphertext[71]                 =   tb_o_ciphertext[70];
assign   tb_o_tag_ready[71]                  =   1'b0;
assign   tb_o_tag[71]                        =   tb_o_tag[70];

// CLK no. 72/1240
// *************************************************
assign   tb_i_valid[72]                      =   1'b0;
assign   tb_i_reset[72]                      =   1'b0;
assign   tb_i_sop[72]                        =   1'b0;
assign   tb_i_key_update[72]                 =   1'b0;
assign   tb_i_key[72]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[72]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[72]               =   1'b0;
assign   tb_i_rf_static_encrypt[72]          =   1'b1;
assign   tb_i_clear_fault_flags[72]          =   1'b0;
assign   tb_i_rf_static_aad_length[72]       =   64'h0000000000000100;
assign   tb_i_aad[72]                        =   tb_i_aad[71];
assign   tb_i_rf_static_plaintext_length[72] =   64'h0000000000000280;
assign   tb_i_plaintext[72]                  =   tb_i_plaintext[71];
assign   tb_o_valid[72]                      =   1'b0;
assign   tb_o_sop[72]                        =   1'b0;
assign   tb_o_ciphertext[72]                 =   tb_o_ciphertext[71];
assign   tb_o_tag_ready[72]                  =   1'b0;
assign   tb_o_tag[72]                        =   tb_o_tag[71];

// CLK no. 73/1240
// *************************************************
assign   tb_i_valid[73]                      =   1'b0;
assign   tb_i_reset[73]                      =   1'b0;
assign   tb_i_sop[73]                        =   1'b0;
assign   tb_i_key_update[73]                 =   1'b0;
assign   tb_i_key[73]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[73]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[73]               =   1'b0;
assign   tb_i_rf_static_encrypt[73]          =   1'b1;
assign   tb_i_clear_fault_flags[73]          =   1'b0;
assign   tb_i_rf_static_aad_length[73]       =   64'h0000000000000100;
assign   tb_i_aad[73]                        =   tb_i_aad[72];
assign   tb_i_rf_static_plaintext_length[73] =   64'h0000000000000280;
assign   tb_i_plaintext[73]                  =   tb_i_plaintext[72];
assign   tb_o_valid[73]                      =   1'b0;
assign   tb_o_sop[73]                        =   1'b0;
assign   tb_o_ciphertext[73]                 =   tb_o_ciphertext[72];
assign   tb_o_tag_ready[73]                  =   1'b0;
assign   tb_o_tag[73]                        =   tb_o_tag[72];

// CLK no. 74/1240
// *************************************************
assign   tb_i_valid[74]                      =   1'b0;
assign   tb_i_reset[74]                      =   1'b0;
assign   tb_i_sop[74]                        =   1'b0;
assign   tb_i_key_update[74]                 =   1'b0;
assign   tb_i_key[74]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[74]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[74]               =   1'b0;
assign   tb_i_rf_static_encrypt[74]          =   1'b1;
assign   tb_i_clear_fault_flags[74]          =   1'b0;
assign   tb_i_rf_static_aad_length[74]       =   64'h0000000000000100;
assign   tb_i_aad[74]                        =   tb_i_aad[73];
assign   tb_i_rf_static_plaintext_length[74] =   64'h0000000000000280;
assign   tb_i_plaintext[74]                  =   tb_i_plaintext[73];
assign   tb_o_valid[74]                      =   1'b0;
assign   tb_o_sop[74]                        =   1'b0;
assign   tb_o_ciphertext[74]                 =   tb_o_ciphertext[73];
assign   tb_o_tag_ready[74]                  =   1'b0;
assign   tb_o_tag[74]                        =   tb_o_tag[73];

// CLK no. 75/1240
// *************************************************
assign   tb_i_valid[75]                      =   1'b0;
assign   tb_i_reset[75]                      =   1'b0;
assign   tb_i_sop[75]                        =   1'b0;
assign   tb_i_key_update[75]                 =   1'b0;
assign   tb_i_key[75]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[75]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[75]               =   1'b0;
assign   tb_i_rf_static_encrypt[75]          =   1'b1;
assign   tb_i_clear_fault_flags[75]          =   1'b0;
assign   tb_i_rf_static_aad_length[75]       =   64'h0000000000000100;
assign   tb_i_aad[75]                        =   tb_i_aad[74];
assign   tb_i_rf_static_plaintext_length[75] =   64'h0000000000000280;
assign   tb_i_plaintext[75]                  =   tb_i_plaintext[74];
assign   tb_o_valid[75]                      =   1'b0;
assign   tb_o_sop[75]                        =   1'b0;
assign   tb_o_ciphertext[75]                 =   tb_o_ciphertext[74];
assign   tb_o_tag_ready[75]                  =   1'b0;
assign   tb_o_tag[75]                        =   tb_o_tag[74];

// CLK no. 76/1240
// *************************************************
assign   tb_i_valid[76]                      =   1'b0;
assign   tb_i_reset[76]                      =   1'b0;
assign   tb_i_sop[76]                        =   1'b0;
assign   tb_i_key_update[76]                 =   1'b0;
assign   tb_i_key[76]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[76]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[76]               =   1'b0;
assign   tb_i_rf_static_encrypt[76]          =   1'b1;
assign   tb_i_clear_fault_flags[76]          =   1'b0;
assign   tb_i_rf_static_aad_length[76]       =   64'h0000000000000100;
assign   tb_i_aad[76]                        =   tb_i_aad[75];
assign   tb_i_rf_static_plaintext_length[76] =   64'h0000000000000280;
assign   tb_i_plaintext[76]                  =   tb_i_plaintext[75];
assign   tb_o_valid[76]                      =   1'b0;
assign   tb_o_sop[76]                        =   1'b0;
assign   tb_o_ciphertext[76]                 =   tb_o_ciphertext[75];
assign   tb_o_tag_ready[76]                  =   1'b0;
assign   tb_o_tag[76]                        =   tb_o_tag[75];

// CLK no. 77/1240
// *************************************************
assign   tb_i_valid[77]                      =   1'b0;
assign   tb_i_reset[77]                      =   1'b0;
assign   tb_i_sop[77]                        =   1'b0;
assign   tb_i_key_update[77]                 =   1'b0;
assign   tb_i_key[77]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[77]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[77]               =   1'b0;
assign   tb_i_rf_static_encrypt[77]          =   1'b1;
assign   tb_i_clear_fault_flags[77]          =   1'b0;
assign   tb_i_rf_static_aad_length[77]       =   64'h0000000000000100;
assign   tb_i_aad[77]                        =   tb_i_aad[76];
assign   tb_i_rf_static_plaintext_length[77] =   64'h0000000000000280;
assign   tb_i_plaintext[77]                  =   tb_i_plaintext[76];
assign   tb_o_valid[77]                      =   1'b0;
assign   tb_o_sop[77]                        =   1'b0;
assign   tb_o_ciphertext[77]                 =   tb_o_ciphertext[76];
assign   tb_o_tag_ready[77]                  =   1'b0;
assign   tb_o_tag[77]                        =   tb_o_tag[76];

// CLK no. 78/1240
// *************************************************
assign   tb_i_valid[78]                      =   1'b0;
assign   tb_i_reset[78]                      =   1'b0;
assign   tb_i_sop[78]                        =   1'b0;
assign   tb_i_key_update[78]                 =   1'b0;
assign   tb_i_key[78]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[78]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[78]               =   1'b0;
assign   tb_i_rf_static_encrypt[78]          =   1'b1;
assign   tb_i_clear_fault_flags[78]          =   1'b0;
assign   tb_i_rf_static_aad_length[78]       =   64'h0000000000000100;
assign   tb_i_aad[78]                        =   tb_i_aad[77];
assign   tb_i_rf_static_plaintext_length[78] =   64'h0000000000000280;
assign   tb_i_plaintext[78]                  =   tb_i_plaintext[77];
assign   tb_o_valid[78]                      =   1'b0;
assign   tb_o_sop[78]                        =   1'b0;
assign   tb_o_ciphertext[78]                 =   tb_o_ciphertext[77];
assign   tb_o_tag_ready[78]                  =   1'b0;
assign   tb_o_tag[78]                        =   tb_o_tag[77];

// CLK no. 79/1240
// *************************************************
assign   tb_i_valid[79]                      =   1'b0;
assign   tb_i_reset[79]                      =   1'b0;
assign   tb_i_sop[79]                        =   1'b0;
assign   tb_i_key_update[79]                 =   1'b0;
assign   tb_i_key[79]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[79]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[79]               =   1'b0;
assign   tb_i_rf_static_encrypt[79]          =   1'b1;
assign   tb_i_clear_fault_flags[79]          =   1'b0;
assign   tb_i_rf_static_aad_length[79]       =   64'h0000000000000100;
assign   tb_i_aad[79]                        =   tb_i_aad[78];
assign   tb_i_rf_static_plaintext_length[79] =   64'h0000000000000280;
assign   tb_i_plaintext[79]                  =   tb_i_plaintext[78];
assign   tb_o_valid[79]                      =   1'b0;
assign   tb_o_sop[79]                        =   1'b0;
assign   tb_o_ciphertext[79]                 =   tb_o_ciphertext[78];
assign   tb_o_tag_ready[79]                  =   1'b0;
assign   tb_o_tag[79]                        =   tb_o_tag[78];

// CLK no. 80/1240
// *************************************************
assign   tb_i_valid[80]                      =   1'b0;
assign   tb_i_reset[80]                      =   1'b0;
assign   tb_i_sop[80]                        =   1'b0;
assign   tb_i_key_update[80]                 =   1'b0;
assign   tb_i_key[80]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[80]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[80]               =   1'b0;
assign   tb_i_rf_static_encrypt[80]          =   1'b1;
assign   tb_i_clear_fault_flags[80]          =   1'b0;
assign   tb_i_rf_static_aad_length[80]       =   64'h0000000000000100;
assign   tb_i_aad[80]                        =   tb_i_aad[79];
assign   tb_i_rf_static_plaintext_length[80] =   64'h0000000000000280;
assign   tb_i_plaintext[80]                  =   tb_i_plaintext[79];
assign   tb_o_valid[80]                      =   1'b0;
assign   tb_o_sop[80]                        =   1'b0;
assign   tb_o_ciphertext[80]                 =   tb_o_ciphertext[79];
assign   tb_o_tag_ready[80]                  =   1'b0;
assign   tb_o_tag[80]                        =   tb_o_tag[79];

// CLK no. 81/1240
// *************************************************
assign   tb_i_valid[81]                      =   1'b0;
assign   tb_i_reset[81]                      =   1'b0;
assign   tb_i_sop[81]                        =   1'b0;
assign   tb_i_key_update[81]                 =   1'b0;
assign   tb_i_key[81]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[81]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[81]               =   1'b0;
assign   tb_i_rf_static_encrypt[81]          =   1'b1;
assign   tb_i_clear_fault_flags[81]          =   1'b0;
assign   tb_i_rf_static_aad_length[81]       =   64'h0000000000000100;
assign   tb_i_aad[81]                        =   tb_i_aad[80];
assign   tb_i_rf_static_plaintext_length[81] =   64'h0000000000000280;
assign   tb_i_plaintext[81]                  =   tb_i_plaintext[80];
assign   tb_o_valid[81]                      =   1'b0;
assign   tb_o_sop[81]                        =   1'b0;
assign   tb_o_ciphertext[81]                 =   tb_o_ciphertext[80];
assign   tb_o_tag_ready[81]                  =   1'b0;
assign   tb_o_tag[81]                        =   tb_o_tag[80];

// CLK no. 82/1240
// *************************************************
assign   tb_i_valid[82]                      =   1'b0;
assign   tb_i_reset[82]                      =   1'b0;
assign   tb_i_sop[82]                        =   1'b0;
assign   tb_i_key_update[82]                 =   1'b0;
assign   tb_i_key[82]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[82]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[82]               =   1'b0;
assign   tb_i_rf_static_encrypt[82]          =   1'b1;
assign   tb_i_clear_fault_flags[82]          =   1'b0;
assign   tb_i_rf_static_aad_length[82]       =   64'h0000000000000100;
assign   tb_i_aad[82]                        =   tb_i_aad[81];
assign   tb_i_rf_static_plaintext_length[82] =   64'h0000000000000280;
assign   tb_i_plaintext[82]                  =   tb_i_plaintext[81];
assign   tb_o_valid[82]                      =   1'b0;
assign   tb_o_sop[82]                        =   1'b0;
assign   tb_o_ciphertext[82]                 =   tb_o_ciphertext[81];
assign   tb_o_tag_ready[82]                  =   1'b0;
assign   tb_o_tag[82]                        =   tb_o_tag[81];

// CLK no. 83/1240
// *************************************************
assign   tb_i_valid[83]                      =   1'b0;
assign   tb_i_reset[83]                      =   1'b0;
assign   tb_i_sop[83]                        =   1'b0;
assign   tb_i_key_update[83]                 =   1'b0;
assign   tb_i_key[83]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[83]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[83]               =   1'b0;
assign   tb_i_rf_static_encrypt[83]          =   1'b1;
assign   tb_i_clear_fault_flags[83]          =   1'b0;
assign   tb_i_rf_static_aad_length[83]       =   64'h0000000000000100;
assign   tb_i_aad[83]                        =   tb_i_aad[82];
assign   tb_i_rf_static_plaintext_length[83] =   64'h0000000000000280;
assign   tb_i_plaintext[83]                  =   tb_i_plaintext[82];
assign   tb_o_valid[83]                      =   1'b0;
assign   tb_o_sop[83]                        =   1'b0;
assign   tb_o_ciphertext[83]                 =   tb_o_ciphertext[82];
assign   tb_o_tag_ready[83]                  =   1'b0;
assign   tb_o_tag[83]                        =   tb_o_tag[82];

// CLK no. 84/1240
// *************************************************
assign   tb_i_valid[84]                      =   1'b0;
assign   tb_i_reset[84]                      =   1'b0;
assign   tb_i_sop[84]                        =   1'b0;
assign   tb_i_key_update[84]                 =   1'b0;
assign   tb_i_key[84]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[84]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[84]               =   1'b0;
assign   tb_i_rf_static_encrypt[84]          =   1'b1;
assign   tb_i_clear_fault_flags[84]          =   1'b0;
assign   tb_i_rf_static_aad_length[84]       =   64'h0000000000000100;
assign   tb_i_aad[84]                        =   tb_i_aad[83];
assign   tb_i_rf_static_plaintext_length[84] =   64'h0000000000000280;
assign   tb_i_plaintext[84]                  =   tb_i_plaintext[83];
assign   tb_o_valid[84]                      =   1'b0;
assign   tb_o_sop[84]                        =   1'b0;
assign   tb_o_ciphertext[84]                 =   tb_o_ciphertext[83];
assign   tb_o_tag_ready[84]                  =   1'b0;
assign   tb_o_tag[84]                        =   tb_o_tag[83];

// CLK no. 85/1240
// *************************************************
assign   tb_i_valid[85]                      =   1'b0;
assign   tb_i_reset[85]                      =   1'b0;
assign   tb_i_sop[85]                        =   1'b0;
assign   tb_i_key_update[85]                 =   1'b0;
assign   tb_i_key[85]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[85]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[85]               =   1'b0;
assign   tb_i_rf_static_encrypt[85]          =   1'b1;
assign   tb_i_clear_fault_flags[85]          =   1'b0;
assign   tb_i_rf_static_aad_length[85]       =   64'h0000000000000100;
assign   tb_i_aad[85]                        =   tb_i_aad[84];
assign   tb_i_rf_static_plaintext_length[85] =   64'h0000000000000280;
assign   tb_i_plaintext[85]                  =   tb_i_plaintext[84];
assign   tb_o_valid[85]                      =   1'b0;
assign   tb_o_sop[85]                        =   1'b0;
assign   tb_o_ciphertext[85]                 =   tb_o_ciphertext[84];
assign   tb_o_tag_ready[85]                  =   1'b0;
assign   tb_o_tag[85]                        =   tb_o_tag[84];

// CLK no. 86/1240
// *************************************************
assign   tb_i_valid[86]                      =   1'b0;
assign   tb_i_reset[86]                      =   1'b0;
assign   tb_i_sop[86]                        =   1'b0;
assign   tb_i_key_update[86]                 =   1'b0;
assign   tb_i_key[86]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[86]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[86]               =   1'b0;
assign   tb_i_rf_static_encrypt[86]          =   1'b1;
assign   tb_i_clear_fault_flags[86]          =   1'b0;
assign   tb_i_rf_static_aad_length[86]       =   64'h0000000000000100;
assign   tb_i_aad[86]                        =   tb_i_aad[85];
assign   tb_i_rf_static_plaintext_length[86] =   64'h0000000000000280;
assign   tb_i_plaintext[86]                  =   tb_i_plaintext[85];
assign   tb_o_valid[86]                      =   1'b0;
assign   tb_o_sop[86]                        =   1'b0;
assign   tb_o_ciphertext[86]                 =   tb_o_ciphertext[85];
assign   tb_o_tag_ready[86]                  =   1'b0;
assign   tb_o_tag[86]                        =   tb_o_tag[85];

// CLK no. 87/1240
// *************************************************
assign   tb_i_valid[87]                      =   1'b0;
assign   tb_i_reset[87]                      =   1'b0;
assign   tb_i_sop[87]                        =   1'b0;
assign   tb_i_key_update[87]                 =   1'b0;
assign   tb_i_key[87]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[87]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[87]               =   1'b0;
assign   tb_i_rf_static_encrypt[87]          =   1'b1;
assign   tb_i_clear_fault_flags[87]          =   1'b0;
assign   tb_i_rf_static_aad_length[87]       =   64'h0000000000000100;
assign   tb_i_aad[87]                        =   tb_i_aad[86];
assign   tb_i_rf_static_plaintext_length[87] =   64'h0000000000000280;
assign   tb_i_plaintext[87]                  =   tb_i_plaintext[86];
assign   tb_o_valid[87]                      =   1'b0;
assign   tb_o_sop[87]                        =   1'b0;
assign   tb_o_ciphertext[87]                 =   tb_o_ciphertext[86];
assign   tb_o_tag_ready[87]                  =   1'b0;
assign   tb_o_tag[87]                        =   tb_o_tag[86];

// CLK no. 88/1240
// *************************************************
assign   tb_i_valid[88]                      =   1'b0;
assign   tb_i_reset[88]                      =   1'b0;
assign   tb_i_sop[88]                        =   1'b0;
assign   tb_i_key_update[88]                 =   1'b0;
assign   tb_i_key[88]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[88]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[88]               =   1'b0;
assign   tb_i_rf_static_encrypt[88]          =   1'b1;
assign   tb_i_clear_fault_flags[88]          =   1'b0;
assign   tb_i_rf_static_aad_length[88]       =   64'h0000000000000100;
assign   tb_i_aad[88]                        =   tb_i_aad[87];
assign   tb_i_rf_static_plaintext_length[88] =   64'h0000000000000280;
assign   tb_i_plaintext[88]                  =   tb_i_plaintext[87];
assign   tb_o_valid[88]                      =   1'b0;
assign   tb_o_sop[88]                        =   1'b0;
assign   tb_o_ciphertext[88]                 =   tb_o_ciphertext[87];
assign   tb_o_tag_ready[88]                  =   1'b0;
assign   tb_o_tag[88]                        =   tb_o_tag[87];

// CLK no. 89/1240
// *************************************************
assign   tb_i_valid[89]                      =   1'b0;
assign   tb_i_reset[89]                      =   1'b0;
assign   tb_i_sop[89]                        =   1'b0;
assign   tb_i_key_update[89]                 =   1'b0;
assign   tb_i_key[89]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[89]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[89]               =   1'b0;
assign   tb_i_rf_static_encrypt[89]          =   1'b1;
assign   tb_i_clear_fault_flags[89]          =   1'b0;
assign   tb_i_rf_static_aad_length[89]       =   64'h0000000000000100;
assign   tb_i_aad[89]                        =   tb_i_aad[88];
assign   tb_i_rf_static_plaintext_length[89] =   64'h0000000000000280;
assign   tb_i_plaintext[89]                  =   tb_i_plaintext[88];
assign   tb_o_valid[89]                      =   1'b0;
assign   tb_o_sop[89]                        =   1'b0;
assign   tb_o_ciphertext[89]                 =   tb_o_ciphertext[88];
assign   tb_o_tag_ready[89]                  =   1'b0;
assign   tb_o_tag[89]                        =   tb_o_tag[88];

// CLK no. 90/1240
// *************************************************
assign   tb_i_valid[90]                      =   1'b0;
assign   tb_i_reset[90]                      =   1'b0;
assign   tb_i_sop[90]                        =   1'b0;
assign   tb_i_key_update[90]                 =   1'b0;
assign   tb_i_key[90]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[90]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[90]               =   1'b0;
assign   tb_i_rf_static_encrypt[90]          =   1'b1;
assign   tb_i_clear_fault_flags[90]          =   1'b0;
assign   tb_i_rf_static_aad_length[90]       =   64'h0000000000000100;
assign   tb_i_aad[90]                        =   tb_i_aad[89];
assign   tb_i_rf_static_plaintext_length[90] =   64'h0000000000000280;
assign   tb_i_plaintext[90]                  =   tb_i_plaintext[89];
assign   tb_o_valid[90]                      =   1'b0;
assign   tb_o_sop[90]                        =   1'b0;
assign   tb_o_ciphertext[90]                 =   tb_o_ciphertext[89];
assign   tb_o_tag_ready[90]                  =   1'b0;
assign   tb_o_tag[90]                        =   tb_o_tag[89];

// CLK no. 91/1240
// *************************************************
assign   tb_i_valid[91]                      =   1'b0;
assign   tb_i_reset[91]                      =   1'b0;
assign   tb_i_sop[91]                        =   1'b0;
assign   tb_i_key_update[91]                 =   1'b0;
assign   tb_i_key[91]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[91]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[91]               =   1'b0;
assign   tb_i_rf_static_encrypt[91]          =   1'b1;
assign   tb_i_clear_fault_flags[91]          =   1'b0;
assign   tb_i_rf_static_aad_length[91]       =   64'h0000000000000100;
assign   tb_i_aad[91]                        =   tb_i_aad[90];
assign   tb_i_rf_static_plaintext_length[91] =   64'h0000000000000280;
assign   tb_i_plaintext[91]                  =   tb_i_plaintext[90];
assign   tb_o_valid[91]                      =   1'b0;
assign   tb_o_sop[91]                        =   1'b0;
assign   tb_o_ciphertext[91]                 =   tb_o_ciphertext[90];
assign   tb_o_tag_ready[91]                  =   1'b0;
assign   tb_o_tag[91]                        =   tb_o_tag[90];

// CLK no. 92/1240
// *************************************************
assign   tb_i_valid[92]                      =   1'b0;
assign   tb_i_reset[92]                      =   1'b0;
assign   tb_i_sop[92]                        =   1'b0;
assign   tb_i_key_update[92]                 =   1'b0;
assign   tb_i_key[92]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[92]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[92]               =   1'b0;
assign   tb_i_rf_static_encrypt[92]          =   1'b1;
assign   tb_i_clear_fault_flags[92]          =   1'b0;
assign   tb_i_rf_static_aad_length[92]       =   64'h0000000000000100;
assign   tb_i_aad[92]                        =   tb_i_aad[91];
assign   tb_i_rf_static_plaintext_length[92] =   64'h0000000000000280;
assign   tb_i_plaintext[92]                  =   tb_i_plaintext[91];
assign   tb_o_valid[92]                      =   1'b0;
assign   tb_o_sop[92]                        =   1'b0;
assign   tb_o_ciphertext[92]                 =   tb_o_ciphertext[91];
assign   tb_o_tag_ready[92]                  =   1'b0;
assign   tb_o_tag[92]                        =   tb_o_tag[91];

// CLK no. 93/1240
// *************************************************
assign   tb_i_valid[93]                      =   1'b0;
assign   tb_i_reset[93]                      =   1'b0;
assign   tb_i_sop[93]                        =   1'b0;
assign   tb_i_key_update[93]                 =   1'b0;
assign   tb_i_key[93]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[93]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[93]               =   1'b0;
assign   tb_i_rf_static_encrypt[93]          =   1'b1;
assign   tb_i_clear_fault_flags[93]          =   1'b0;
assign   tb_i_rf_static_aad_length[93]       =   64'h0000000000000100;
assign   tb_i_aad[93]                        =   tb_i_aad[92];
assign   tb_i_rf_static_plaintext_length[93] =   64'h0000000000000280;
assign   tb_i_plaintext[93]                  =   tb_i_plaintext[92];
assign   tb_o_valid[93]                      =   1'b0;
assign   tb_o_sop[93]                        =   1'b0;
assign   tb_o_ciphertext[93]                 =   tb_o_ciphertext[92];
assign   tb_o_tag_ready[93]                  =   1'b0;
assign   tb_o_tag[93]                        =   tb_o_tag[92];

// CLK no. 94/1240
// *************************************************
assign   tb_i_valid[94]                      =   1'b0;
assign   tb_i_reset[94]                      =   1'b0;
assign   tb_i_sop[94]                        =   1'b0;
assign   tb_i_key_update[94]                 =   1'b0;
assign   tb_i_key[94]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[94]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[94]               =   1'b0;
assign   tb_i_rf_static_encrypt[94]          =   1'b1;
assign   tb_i_clear_fault_flags[94]          =   1'b0;
assign   tb_i_rf_static_aad_length[94]       =   64'h0000000000000100;
assign   tb_i_aad[94]                        =   tb_i_aad[93];
assign   tb_i_rf_static_plaintext_length[94] =   64'h0000000000000280;
assign   tb_i_plaintext[94]                  =   tb_i_plaintext[93];
assign   tb_o_valid[94]                      =   1'b0;
assign   tb_o_sop[94]                        =   1'b0;
assign   tb_o_ciphertext[94]                 =   tb_o_ciphertext[93];
assign   tb_o_tag_ready[94]                  =   1'b0;
assign   tb_o_tag[94]                        =   tb_o_tag[93];

// CLK no. 95/1240
// *************************************************
assign   tb_i_valid[95]                      =   1'b0;
assign   tb_i_reset[95]                      =   1'b0;
assign   tb_i_sop[95]                        =   1'b0;
assign   tb_i_key_update[95]                 =   1'b0;
assign   tb_i_key[95]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[95]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[95]               =   1'b0;
assign   tb_i_rf_static_encrypt[95]          =   1'b1;
assign   tb_i_clear_fault_flags[95]          =   1'b0;
assign   tb_i_rf_static_aad_length[95]       =   64'h0000000000000100;
assign   tb_i_aad[95]                        =   tb_i_aad[94];
assign   tb_i_rf_static_plaintext_length[95] =   64'h0000000000000280;
assign   tb_i_plaintext[95]                  =   tb_i_plaintext[94];
assign   tb_o_valid[95]                      =   1'b0;
assign   tb_o_sop[95]                        =   1'b0;
assign   tb_o_ciphertext[95]                 =   tb_o_ciphertext[94];
assign   tb_o_tag_ready[95]                  =   1'b0;
assign   tb_o_tag[95]                        =   tb_o_tag[94];

// CLK no. 96/1240
// *************************************************
assign   tb_i_valid[96]                      =   1'b0;
assign   tb_i_reset[96]                      =   1'b0;
assign   tb_i_sop[96]                        =   1'b0;
assign   tb_i_key_update[96]                 =   1'b0;
assign   tb_i_key[96]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[96]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[96]               =   1'b0;
assign   tb_i_rf_static_encrypt[96]          =   1'b1;
assign   tb_i_clear_fault_flags[96]          =   1'b0;
assign   tb_i_rf_static_aad_length[96]       =   64'h0000000000000100;
assign   tb_i_aad[96]                        =   tb_i_aad[95];
assign   tb_i_rf_static_plaintext_length[96] =   64'h0000000000000280;
assign   tb_i_plaintext[96]                  =   tb_i_plaintext[95];
assign   tb_o_valid[96]                      =   1'b0;
assign   tb_o_sop[96]                        =   1'b0;
assign   tb_o_ciphertext[96]                 =   tb_o_ciphertext[95];
assign   tb_o_tag_ready[96]                  =   1'b0;
assign   tb_o_tag[96]                        =   tb_o_tag[95];

// CLK no. 97/1240
// *************************************************
assign   tb_i_valid[97]                      =   1'b0;
assign   tb_i_reset[97]                      =   1'b0;
assign   tb_i_sop[97]                        =   1'b0;
assign   tb_i_key_update[97]                 =   1'b0;
assign   tb_i_key[97]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[97]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[97]               =   1'b0;
assign   tb_i_rf_static_encrypt[97]          =   1'b1;
assign   tb_i_clear_fault_flags[97]          =   1'b0;
assign   tb_i_rf_static_aad_length[97]       =   64'h0000000000000100;
assign   tb_i_aad[97]                        =   tb_i_aad[96];
assign   tb_i_rf_static_plaintext_length[97] =   64'h0000000000000280;
assign   tb_i_plaintext[97]                  =   tb_i_plaintext[96];
assign   tb_o_valid[97]                      =   1'b0;
assign   tb_o_sop[97]                        =   1'b0;
assign   tb_o_ciphertext[97]                 =   tb_o_ciphertext[96];
assign   tb_o_tag_ready[97]                  =   1'b0;
assign   tb_o_tag[97]                        =   tb_o_tag[96];

// CLK no. 98/1240
// *************************************************
assign   tb_i_valid[98]                      =   1'b0;
assign   tb_i_reset[98]                      =   1'b0;
assign   tb_i_sop[98]                        =   1'b0;
assign   tb_i_key_update[98]                 =   1'b0;
assign   tb_i_key[98]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[98]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[98]               =   1'b0;
assign   tb_i_rf_static_encrypt[98]          =   1'b1;
assign   tb_i_clear_fault_flags[98]          =   1'b0;
assign   tb_i_rf_static_aad_length[98]       =   64'h0000000000000100;
assign   tb_i_aad[98]                        =   tb_i_aad[97];
assign   tb_i_rf_static_plaintext_length[98] =   64'h0000000000000280;
assign   tb_i_plaintext[98]                  =   tb_i_plaintext[97];
assign   tb_o_valid[98]                      =   1'b0;
assign   tb_o_sop[98]                        =   1'b0;
assign   tb_o_ciphertext[98]                 =   tb_o_ciphertext[97];
assign   tb_o_tag_ready[98]                  =   1'b0;
assign   tb_o_tag[98]                        =   tb_o_tag[97];

// CLK no. 99/1240
// *************************************************
assign   tb_i_valid[99]                      =   1'b0;
assign   tb_i_reset[99]                      =   1'b0;
assign   tb_i_sop[99]                        =   1'b0;
assign   tb_i_key_update[99]                 =   1'b0;
assign   tb_i_key[99]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[99]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[99]               =   1'b0;
assign   tb_i_rf_static_encrypt[99]          =   1'b1;
assign   tb_i_clear_fault_flags[99]          =   1'b0;
assign   tb_i_rf_static_aad_length[99]       =   64'h0000000000000100;
assign   tb_i_aad[99]                        =   tb_i_aad[98];
assign   tb_i_rf_static_plaintext_length[99] =   64'h0000000000000280;
assign   tb_i_plaintext[99]                  =   tb_i_plaintext[98];
assign   tb_o_valid[99]                      =   1'b0;
assign   tb_o_sop[99]                        =   1'b0;
assign   tb_o_ciphertext[99]                 =   tb_o_ciphertext[98];
assign   tb_o_tag_ready[99]                  =   1'b0;
assign   tb_o_tag[99]                        =   tb_o_tag[98];

// CLK no. 100/1240
// *************************************************
assign   tb_i_valid[100]                      =   1'b0;
assign   tb_i_reset[100]                      =   1'b0;
assign   tb_i_sop[100]                        =   1'b0;
assign   tb_i_key_update[100]                 =   1'b0;
assign   tb_i_key[100]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[100]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[100]               =   1'b0;
assign   tb_i_rf_static_encrypt[100]          =   1'b1;
assign   tb_i_clear_fault_flags[100]          =   1'b0;
assign   tb_i_rf_static_aad_length[100]       =   64'h0000000000000100;
assign   tb_i_aad[100]                        =   tb_i_aad[99];
assign   tb_i_rf_static_plaintext_length[100] =   64'h0000000000000280;
assign   tb_i_plaintext[100]                  =   tb_i_plaintext[99];
assign   tb_o_valid[100]                      =   1'b0;
assign   tb_o_sop[100]                        =   1'b0;
assign   tb_o_ciphertext[100]                 =   tb_o_ciphertext[99];
assign   tb_o_tag_ready[100]                  =   1'b0;
assign   tb_o_tag[100]                        =   tb_o_tag[99];

// CLK no. 101/1240
// *************************************************
assign   tb_i_valid[101]                      =   1'b0;
assign   tb_i_reset[101]                      =   1'b0;
assign   tb_i_sop[101]                        =   1'b0;
assign   tb_i_key_update[101]                 =   1'b0;
assign   tb_i_key[101]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[101]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[101]               =   1'b0;
assign   tb_i_rf_static_encrypt[101]          =   1'b1;
assign   tb_i_clear_fault_flags[101]          =   1'b0;
assign   tb_i_rf_static_aad_length[101]       =   64'h0000000000000100;
assign   tb_i_aad[101]                        =   tb_i_aad[100];
assign   tb_i_rf_static_plaintext_length[101] =   64'h0000000000000280;
assign   tb_i_plaintext[101]                  =   tb_i_plaintext[100];
assign   tb_o_valid[101]                      =   1'b0;
assign   tb_o_sop[101]                        =   1'b0;
assign   tb_o_ciphertext[101]                 =   tb_o_ciphertext[100];
assign   tb_o_tag_ready[101]                  =   1'b0;
assign   tb_o_tag[101]                        =   tb_o_tag[100];

// CLK no. 102/1240
// *************************************************
assign   tb_i_valid[102]                      =   1'b0;
assign   tb_i_reset[102]                      =   1'b0;
assign   tb_i_sop[102]                        =   1'b0;
assign   tb_i_key_update[102]                 =   1'b0;
assign   tb_i_key[102]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[102]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[102]               =   1'b0;
assign   tb_i_rf_static_encrypt[102]          =   1'b1;
assign   tb_i_clear_fault_flags[102]          =   1'b0;
assign   tb_i_rf_static_aad_length[102]       =   64'h0000000000000100;
assign   tb_i_aad[102]                        =   tb_i_aad[101];
assign   tb_i_rf_static_plaintext_length[102] =   64'h0000000000000280;
assign   tb_i_plaintext[102]                  =   tb_i_plaintext[101];
assign   tb_o_valid[102]                      =   1'b0;
assign   tb_o_sop[102]                        =   1'b0;
assign   tb_o_ciphertext[102]                 =   tb_o_ciphertext[101];
assign   tb_o_tag_ready[102]                  =   1'b0;
assign   tb_o_tag[102]                        =   tb_o_tag[101];

// CLK no. 103/1240
// *************************************************
assign   tb_i_valid[103]                      =   1'b0;
assign   tb_i_reset[103]                      =   1'b0;
assign   tb_i_sop[103]                        =   1'b0;
assign   tb_i_key_update[103]                 =   1'b0;
assign   tb_i_key[103]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[103]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[103]               =   1'b0;
assign   tb_i_rf_static_encrypt[103]          =   1'b1;
assign   tb_i_clear_fault_flags[103]          =   1'b0;
assign   tb_i_rf_static_aad_length[103]       =   64'h0000000000000100;
assign   tb_i_aad[103]                        =   tb_i_aad[102];
assign   tb_i_rf_static_plaintext_length[103] =   64'h0000000000000280;
assign   tb_i_plaintext[103]                  =   tb_i_plaintext[102];
assign   tb_o_valid[103]                      =   1'b0;
assign   tb_o_sop[103]                        =   1'b0;
assign   tb_o_ciphertext[103]                 =   tb_o_ciphertext[102];
assign   tb_o_tag_ready[103]                  =   1'b0;
assign   tb_o_tag[103]                        =   tb_o_tag[102];

// CLK no. 104/1240
// *************************************************
assign   tb_i_valid[104]                      =   1'b0;
assign   tb_i_reset[104]                      =   1'b0;
assign   tb_i_sop[104]                        =   1'b0;
assign   tb_i_key_update[104]                 =   1'b0;
assign   tb_i_key[104]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[104]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[104]               =   1'b0;
assign   tb_i_rf_static_encrypt[104]          =   1'b1;
assign   tb_i_clear_fault_flags[104]          =   1'b0;
assign   tb_i_rf_static_aad_length[104]       =   64'h0000000000000100;
assign   tb_i_aad[104]                        =   tb_i_aad[103];
assign   tb_i_rf_static_plaintext_length[104] =   64'h0000000000000280;
assign   tb_i_plaintext[104]                  =   tb_i_plaintext[103];
assign   tb_o_valid[104]                      =   1'b0;
assign   tb_o_sop[104]                        =   1'b0;
assign   tb_o_ciphertext[104]                 =   tb_o_ciphertext[103];
assign   tb_o_tag_ready[104]                  =   1'b0;
assign   tb_o_tag[104]                        =   tb_o_tag[103];

// CLK no. 105/1240
// *************************************************
assign   tb_i_valid[105]                      =   1'b0;
assign   tb_i_reset[105]                      =   1'b0;
assign   tb_i_sop[105]                        =   1'b0;
assign   tb_i_key_update[105]                 =   1'b0;
assign   tb_i_key[105]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[105]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[105]               =   1'b0;
assign   tb_i_rf_static_encrypt[105]          =   1'b1;
assign   tb_i_clear_fault_flags[105]          =   1'b0;
assign   tb_i_rf_static_aad_length[105]       =   64'h0000000000000100;
assign   tb_i_aad[105]                        =   tb_i_aad[104];
assign   tb_i_rf_static_plaintext_length[105] =   64'h0000000000000280;
assign   tb_i_plaintext[105]                  =   tb_i_plaintext[104];
assign   tb_o_valid[105]                      =   1'b0;
assign   tb_o_sop[105]                        =   1'b0;
assign   tb_o_ciphertext[105]                 =   tb_o_ciphertext[104];
assign   tb_o_tag_ready[105]                  =   1'b0;
assign   tb_o_tag[105]                        =   tb_o_tag[104];

// CLK no. 106/1240
// *************************************************
assign   tb_i_valid[106]                      =   1'b0;
assign   tb_i_reset[106]                      =   1'b0;
assign   tb_i_sop[106]                        =   1'b0;
assign   tb_i_key_update[106]                 =   1'b0;
assign   tb_i_key[106]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[106]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[106]               =   1'b0;
assign   tb_i_rf_static_encrypt[106]          =   1'b1;
assign   tb_i_clear_fault_flags[106]          =   1'b0;
assign   tb_i_rf_static_aad_length[106]       =   64'h0000000000000100;
assign   tb_i_aad[106]                        =   tb_i_aad[105];
assign   tb_i_rf_static_plaintext_length[106] =   64'h0000000000000280;
assign   tb_i_plaintext[106]                  =   tb_i_plaintext[105];
assign   tb_o_valid[106]                      =   1'b1;
assign   tb_o_sop[106]                        =   1'b1;
assign   tb_o_ciphertext[106]                 =   256'h3d3778bd93aaf83dac83e8767cc43cda10ff9c7dbfabcdc3e7d89c62655f7bb6;
assign   tb_o_tag_ready[106]                  =   1'b0;
assign   tb_o_tag[106]                        =   tb_o_tag[105];

// CLK no. 107/1240
// *************************************************
assign   tb_i_valid[107]                      =   1'b0;
assign   tb_i_reset[107]                      =   1'b0;
assign   tb_i_sop[107]                        =   1'b0;
assign   tb_i_key_update[107]                 =   1'b0;
assign   tb_i_key[107]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[107]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[107]               =   1'b0;
assign   tb_i_rf_static_encrypt[107]          =   1'b1;
assign   tb_i_clear_fault_flags[107]          =   1'b0;
assign   tb_i_rf_static_aad_length[107]       =   64'h0000000000000100;
assign   tb_i_aad[107]                        =   tb_i_aad[106];
assign   tb_i_rf_static_plaintext_length[107] =   64'h0000000000000280;
assign   tb_i_plaintext[107]                  =   tb_i_plaintext[106];
assign   tb_o_valid[107]                      =   1'b1;
assign   tb_o_sop[107]                        =   1'b0;
assign   tb_o_ciphertext[107]                 =   256'habe55dbe62e9005828cc2bd665f1570773f44816682889e19f4cda071b52533e;
assign   tb_o_tag_ready[107]                  =   1'b0;
assign   tb_o_tag[107]                        =   tb_o_tag[106];

// CLK no. 108/1240
// *************************************************
assign   tb_i_valid[108]                      =   1'b0;
assign   tb_i_reset[108]                      =   1'b0;
assign   tb_i_sop[108]                        =   1'b0;
assign   tb_i_key_update[108]                 =   1'b0;
assign   tb_i_key[108]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[108]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[108]               =   1'b0;
assign   tb_i_rf_static_encrypt[108]          =   1'b1;
assign   tb_i_clear_fault_flags[108]          =   1'b0;
assign   tb_i_rf_static_aad_length[108]       =   64'h0000000000000100;
assign   tb_i_aad[108]                        =   tb_i_aad[107];
assign   tb_i_rf_static_plaintext_length[108] =   64'h0000000000000280;
assign   tb_i_plaintext[108]                  =   tb_i_plaintext[107];
assign   tb_o_valid[108]                      =   1'b1;
assign   tb_o_sop[108]                        =   1'b0;
assign   tb_o_ciphertext[108]                 =   256'h1c24392f2fb2e7bdc76c88d7e9c9cd94;
assign   tb_o_tag_ready[108]                  =   1'b0;
assign   tb_o_tag[108]                        =   tb_o_tag[107];

// CLK no. 109/1240
// *************************************************
assign   tb_i_valid[109]                      =   1'b0;
assign   tb_i_reset[109]                      =   1'b0;
assign   tb_i_sop[109]                        =   1'b0;
assign   tb_i_key_update[109]                 =   1'b0;
assign   tb_i_key[109]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[109]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[109]               =   1'b0;
assign   tb_i_rf_static_encrypt[109]          =   1'b1;
assign   tb_i_clear_fault_flags[109]          =   1'b0;
assign   tb_i_rf_static_aad_length[109]       =   64'h0000000000000100;
assign   tb_i_aad[109]                        =   tb_i_aad[108];
assign   tb_i_rf_static_plaintext_length[109] =   64'h0000000000000280;
assign   tb_i_plaintext[109]                  =   tb_i_plaintext[108];
assign   tb_o_valid[109]                      =   1'b0;
assign   tb_o_sop[109]                        =   1'b0;
assign   tb_o_ciphertext[109]                 =   tb_o_ciphertext[108];
assign   tb_o_tag_ready[109]                  =   1'b0;
assign   tb_o_tag[109]                        =   tb_o_tag[108];

// CLK no. 110/1240
// *************************************************
assign   tb_i_valid[110]                      =   1'b0;
assign   tb_i_reset[110]                      =   1'b0;
assign   tb_i_sop[110]                        =   1'b0;
assign   tb_i_key_update[110]                 =   1'b0;
assign   tb_i_key[110]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[110]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[110]               =   1'b0;
assign   tb_i_rf_static_encrypt[110]          =   1'b1;
assign   tb_i_clear_fault_flags[110]          =   1'b0;
assign   tb_i_rf_static_aad_length[110]       =   64'h0000000000000100;
assign   tb_i_aad[110]                        =   tb_i_aad[109];
assign   tb_i_rf_static_plaintext_length[110] =   64'h0000000000000280;
assign   tb_i_plaintext[110]                  =   tb_i_plaintext[109];
assign   tb_o_valid[110]                      =   1'b0;
assign   tb_o_sop[110]                        =   1'b0;
assign   tb_o_ciphertext[110]                 =   tb_o_ciphertext[109];
assign   tb_o_tag_ready[110]                  =   1'b0;
assign   tb_o_tag[110]                        =   tb_o_tag[109];

// CLK no. 111/1240
// *************************************************
assign   tb_i_valid[111]                      =   1'b0;
assign   tb_i_reset[111]                      =   1'b0;
assign   tb_i_sop[111]                        =   1'b0;
assign   tb_i_key_update[111]                 =   1'b0;
assign   tb_i_key[111]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[111]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[111]               =   1'b0;
assign   tb_i_rf_static_encrypt[111]          =   1'b1;
assign   tb_i_clear_fault_flags[111]          =   1'b0;
assign   tb_i_rf_static_aad_length[111]       =   64'h0000000000000100;
assign   tb_i_aad[111]                        =   tb_i_aad[110];
assign   tb_i_rf_static_plaintext_length[111] =   64'h0000000000000280;
assign   tb_i_plaintext[111]                  =   tb_i_plaintext[110];
assign   tb_o_valid[111]                      =   1'b0;
assign   tb_o_sop[111]                        =   1'b0;
assign   tb_o_ciphertext[111]                 =   tb_o_ciphertext[110];
assign   tb_o_tag_ready[111]                  =   1'b0;
assign   tb_o_tag[111]                        =   tb_o_tag[110];

// CLK no. 112/1240
// *************************************************
assign   tb_i_valid[112]                      =   1'b0;
assign   tb_i_reset[112]                      =   1'b0;
assign   tb_i_sop[112]                        =   1'b0;
assign   tb_i_key_update[112]                 =   1'b0;
assign   tb_i_key[112]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[112]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[112]               =   1'b0;
assign   tb_i_rf_static_encrypt[112]          =   1'b1;
assign   tb_i_clear_fault_flags[112]          =   1'b0;
assign   tb_i_rf_static_aad_length[112]       =   64'h0000000000000100;
assign   tb_i_aad[112]                        =   tb_i_aad[111];
assign   tb_i_rf_static_plaintext_length[112] =   64'h0000000000000280;
assign   tb_i_plaintext[112]                  =   tb_i_plaintext[111];
assign   tb_o_valid[112]                      =   1'b0;
assign   tb_o_sop[112]                        =   1'b0;
assign   tb_o_ciphertext[112]                 =   tb_o_ciphertext[111];
assign   tb_o_tag_ready[112]                  =   1'b0;
assign   tb_o_tag[112]                        =   tb_o_tag[111];

// CLK no. 113/1240
// *************************************************
assign   tb_i_valid[113]                      =   1'b0;
assign   tb_i_reset[113]                      =   1'b0;
assign   tb_i_sop[113]                        =   1'b0;
assign   tb_i_key_update[113]                 =   1'b0;
assign   tb_i_key[113]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[113]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[113]               =   1'b0;
assign   tb_i_rf_static_encrypt[113]          =   1'b1;
assign   tb_i_clear_fault_flags[113]          =   1'b0;
assign   tb_i_rf_static_aad_length[113]       =   64'h0000000000000100;
assign   tb_i_aad[113]                        =   tb_i_aad[112];
assign   tb_i_rf_static_plaintext_length[113] =   64'h0000000000000280;
assign   tb_i_plaintext[113]                  =   tb_i_plaintext[112];
assign   tb_o_valid[113]                      =   1'b0;
assign   tb_o_sop[113]                        =   1'b0;
assign   tb_o_ciphertext[113]                 =   tb_o_ciphertext[112];
assign   tb_o_tag_ready[113]                  =   1'b0;
assign   tb_o_tag[113]                        =   tb_o_tag[112];

// CLK no. 114/1240
// *************************************************
assign   tb_i_valid[114]                      =   1'b0;
assign   tb_i_reset[114]                      =   1'b0;
assign   tb_i_sop[114]                        =   1'b0;
assign   tb_i_key_update[114]                 =   1'b0;
assign   tb_i_key[114]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[114]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[114]               =   1'b0;
assign   tb_i_rf_static_encrypt[114]          =   1'b1;
assign   tb_i_clear_fault_flags[114]          =   1'b0;
assign   tb_i_rf_static_aad_length[114]       =   64'h0000000000000100;
assign   tb_i_aad[114]                        =   tb_i_aad[113];
assign   tb_i_rf_static_plaintext_length[114] =   64'h0000000000000280;
assign   tb_i_plaintext[114]                  =   tb_i_plaintext[113];
assign   tb_o_valid[114]                      =   1'b0;
assign   tb_o_sop[114]                        =   1'b0;
assign   tb_o_ciphertext[114]                 =   tb_o_ciphertext[113];
assign   tb_o_tag_ready[114]                  =   1'b0;
assign   tb_o_tag[114]                        =   tb_o_tag[113];

// CLK no. 115/1240
// *************************************************
assign   tb_i_valid[115]                      =   1'b0;
assign   tb_i_reset[115]                      =   1'b0;
assign   tb_i_sop[115]                        =   1'b0;
assign   tb_i_key_update[115]                 =   1'b0;
assign   tb_i_key[115]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[115]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[115]               =   1'b0;
assign   tb_i_rf_static_encrypt[115]          =   1'b1;
assign   tb_i_clear_fault_flags[115]          =   1'b0;
assign   tb_i_rf_static_aad_length[115]       =   64'h0000000000000100;
assign   tb_i_aad[115]                        =   tb_i_aad[114];
assign   tb_i_rf_static_plaintext_length[115] =   64'h0000000000000280;
assign   tb_i_plaintext[115]                  =   tb_i_plaintext[114];
assign   tb_o_valid[115]                      =   1'b0;
assign   tb_o_sop[115]                        =   1'b0;
assign   tb_o_ciphertext[115]                 =   tb_o_ciphertext[114];
assign   tb_o_tag_ready[115]                  =   1'b0;
assign   tb_o_tag[115]                        =   tb_o_tag[114];

// CLK no. 116/1240
// *************************************************
assign   tb_i_valid[116]                      =   1'b0;
assign   tb_i_reset[116]                      =   1'b0;
assign   tb_i_sop[116]                        =   1'b0;
assign   tb_i_key_update[116]                 =   1'b0;
assign   tb_i_key[116]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[116]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[116]               =   1'b0;
assign   tb_i_rf_static_encrypt[116]          =   1'b1;
assign   tb_i_clear_fault_flags[116]          =   1'b0;
assign   tb_i_rf_static_aad_length[116]       =   64'h0000000000000100;
assign   tb_i_aad[116]                        =   tb_i_aad[115];
assign   tb_i_rf_static_plaintext_length[116] =   64'h0000000000000280;
assign   tb_i_plaintext[116]                  =   tb_i_plaintext[115];
assign   tb_o_valid[116]                      =   1'b0;
assign   tb_o_sop[116]                        =   1'b0;
assign   tb_o_ciphertext[116]                 =   tb_o_ciphertext[115];
assign   tb_o_tag_ready[116]                  =   1'b1;
assign   tb_o_tag[116]                        =   128'h3d336f7edbfefbec557a733c74504efe;

// CLK no. 117/1240
// *************************************************
assign   tb_i_valid[117]                      =   1'b0;
assign   tb_i_reset[117]                      =   1'b0;
assign   tb_i_sop[117]                        =   1'b0;
assign   tb_i_key_update[117]                 =   1'b0;
assign   tb_i_key[117]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[117]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[117]               =   1'b0;
assign   tb_i_rf_static_encrypt[117]          =   1'b1;
assign   tb_i_clear_fault_flags[117]          =   1'b0;
assign   tb_i_rf_static_aad_length[117]       =   64'h0000000000000100;
assign   tb_i_aad[117]                        =   tb_i_aad[116];
assign   tb_i_rf_static_plaintext_length[117] =   64'h0000000000000280;
assign   tb_i_plaintext[117]                  =   tb_i_plaintext[116];
assign   tb_o_valid[117]                      =   1'b0;
assign   tb_o_sop[117]                        =   1'b0;
assign   tb_o_ciphertext[117]                 =   tb_o_ciphertext[116];
assign   tb_o_tag_ready[117]                  =   1'b0;
assign   tb_o_tag[117]                        =   tb_o_tag[116];

// CLK no. 118/1240
// *************************************************
assign   tb_i_valid[118]                      =   1'b0;
assign   tb_i_reset[118]                      =   1'b0;
assign   tb_i_sop[118]                        =   1'b0;
assign   tb_i_key_update[118]                 =   1'b0;
assign   tb_i_key[118]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[118]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[118]               =   1'b0;
assign   tb_i_rf_static_encrypt[118]          =   1'b1;
assign   tb_i_clear_fault_flags[118]          =   1'b0;
assign   tb_i_rf_static_aad_length[118]       =   64'h0000000000000100;
assign   tb_i_aad[118]                        =   tb_i_aad[117];
assign   tb_i_rf_static_plaintext_length[118] =   64'h0000000000000280;
assign   tb_i_plaintext[118]                  =   tb_i_plaintext[117];
assign   tb_o_valid[118]                      =   1'b0;
assign   tb_o_sop[118]                        =   1'b0;
assign   tb_o_ciphertext[118]                 =   tb_o_ciphertext[117];
assign   tb_o_tag_ready[118]                  =   1'b0;
assign   tb_o_tag[118]                        =   tb_o_tag[117];

// CLK no. 119/1240
// *************************************************
assign   tb_i_valid[119]                      =   1'b0;
assign   tb_i_reset[119]                      =   1'b0;
assign   tb_i_sop[119]                        =   1'b1;
assign   tb_i_key_update[119]                 =   1'b0;
assign   tb_i_key[119]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[119]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[119]               =   1'b0;
assign   tb_i_rf_static_encrypt[119]          =   1'b1;
assign   tb_i_clear_fault_flags[119]          =   1'b0;
assign   tb_i_rf_static_aad_length[119]       =   64'h0000000000000100;
assign   tb_i_aad[119]                        =   tb_i_aad[118];
assign   tb_i_rf_static_plaintext_length[119] =   64'h0000000000000280;
assign   tb_i_plaintext[119]                  =   tb_i_plaintext[118];
assign   tb_o_valid[119]                      =   1'b0;
assign   tb_o_sop[119]                        =   1'b0;
assign   tb_o_ciphertext[119]                 =   tb_o_ciphertext[118];
assign   tb_o_tag_ready[119]                  =   1'b0;
assign   tb_o_tag[119]                        =   tb_o_tag[118];

// CLK no. 120/1240
// *************************************************
assign   tb_i_valid[120]                      =   1'b1;
assign   tb_i_reset[120]                      =   1'b0;
assign   tb_i_sop[120]                        =   1'b0;
assign   tb_i_key_update[120]                 =   1'b0;
assign   tb_i_key[120]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[120]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[120]               =   1'b0;
assign   tb_i_rf_static_encrypt[120]          =   1'b1;
assign   tb_i_clear_fault_flags[120]          =   1'b0;
assign   tb_i_rf_static_aad_length[120]       =   64'h0000000000000100;
assign   tb_i_aad[120]                        =   256'h474faf91e07f7e6a36d88ba80f126211ec7198b4e7fe60824e2b993af955a1ba;
assign   tb_i_rf_static_plaintext_length[120] =   64'h0000000000000280;
assign   tb_i_plaintext[120]                  =   tb_i_plaintext[119];
assign   tb_o_valid[120]                      =   1'b0;
assign   tb_o_sop[120]                        =   1'b0;
assign   tb_o_ciphertext[120]                 =   tb_o_ciphertext[119];
assign   tb_o_tag_ready[120]                  =   1'b0;
assign   tb_o_tag[120]                        =   tb_o_tag[119];

// CLK no. 121/1240
// *************************************************
assign   tb_i_valid[121]                      =   1'b1;
assign   tb_i_reset[121]                      =   1'b0;
assign   tb_i_sop[121]                        =   1'b0;
assign   tb_i_key_update[121]                 =   1'b0;
assign   tb_i_key[121]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[121]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[121]               =   1'b0;
assign   tb_i_rf_static_encrypt[121]          =   1'b1;
assign   tb_i_clear_fault_flags[121]          =   1'b0;
assign   tb_i_rf_static_aad_length[121]       =   64'h0000000000000100;
assign   tb_i_aad[121]                        =   tb_i_aad[120];
assign   tb_i_rf_static_plaintext_length[121] =   64'h0000000000000280;
assign   tb_i_plaintext[121]                  =   256'h8b5a97fc4a24e77dff1c1a8dac621d59f24706e2a2c67099a226c1cebca3810f;
assign   tb_o_valid[121]                      =   1'b0;
assign   tb_o_sop[121]                        =   1'b0;
assign   tb_o_ciphertext[121]                 =   tb_o_ciphertext[120];
assign   tb_o_tag_ready[121]                  =   1'b0;
assign   tb_o_tag[121]                        =   tb_o_tag[120];

// CLK no. 122/1240
// *************************************************
assign   tb_i_valid[122]                      =   1'b1;
assign   tb_i_reset[122]                      =   1'b0;
assign   tb_i_sop[122]                        =   1'b0;
assign   tb_i_key_update[122]                 =   1'b0;
assign   tb_i_key[122]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[122]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[122]               =   1'b0;
assign   tb_i_rf_static_encrypt[122]          =   1'b1;
assign   tb_i_clear_fault_flags[122]          =   1'b0;
assign   tb_i_rf_static_aad_length[122]       =   64'h0000000000000100;
assign   tb_i_aad[122]                        =   tb_i_aad[121];
assign   tb_i_rf_static_plaintext_length[122] =   64'h0000000000000280;
assign   tb_i_plaintext[122]                  =   256'h2d5a278ee0443011bbdf6ec0b6d147c4c0e8eb0c93fe17c756d1dfdb18788d25;
assign   tb_o_valid[122]                      =   1'b0;
assign   tb_o_sop[122]                        =   1'b0;
assign   tb_o_ciphertext[122]                 =   tb_o_ciphertext[121];
assign   tb_o_tag_ready[122]                  =   1'b0;
assign   tb_o_tag[122]                        =   tb_o_tag[121];

// CLK no. 123/1240
// *************************************************
assign   tb_i_valid[123]                      =   1'b1;
assign   tb_i_reset[123]                      =   1'b0;
assign   tb_i_sop[123]                        =   1'b0;
assign   tb_i_key_update[123]                 =   1'b0;
assign   tb_i_key[123]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[123]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[123]               =   1'b0;
assign   tb_i_rf_static_encrypt[123]          =   1'b1;
assign   tb_i_clear_fault_flags[123]          =   1'b0;
assign   tb_i_rf_static_aad_length[123]       =   64'h0000000000000100;
assign   tb_i_aad[123]                        =   tb_i_aad[122];
assign   tb_i_rf_static_plaintext_length[123] =   64'h0000000000000280;
assign   tb_i_plaintext[123]                  =   256'he440b42d629532fc46bb38bc46756bff;
assign   tb_o_valid[123]                      =   1'b0;
assign   tb_o_sop[123]                        =   1'b0;
assign   tb_o_ciphertext[123]                 =   tb_o_ciphertext[122];
assign   tb_o_tag_ready[123]                  =   1'b0;
assign   tb_o_tag[123]                        =   tb_o_tag[122];

// CLK no. 124/1240
// *************************************************
assign   tb_i_valid[124]                      =   1'b0;
assign   tb_i_reset[124]                      =   1'b0;
assign   tb_i_sop[124]                        =   1'b0;
assign   tb_i_key_update[124]                 =   1'b0;
assign   tb_i_key[124]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[124]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[124]               =   1'b0;
assign   tb_i_rf_static_encrypt[124]          =   1'b1;
assign   tb_i_clear_fault_flags[124]          =   1'b0;
assign   tb_i_rf_static_aad_length[124]       =   64'h0000000000000100;
assign   tb_i_aad[124]                        =   tb_i_aad[123];
assign   tb_i_rf_static_plaintext_length[124] =   64'h0000000000000280;
assign   tb_i_plaintext[124]                  =   tb_i_plaintext[123];
assign   tb_o_valid[124]                      =   1'b0;
assign   tb_o_sop[124]                        =   1'b0;
assign   tb_o_ciphertext[124]                 =   tb_o_ciphertext[123];
assign   tb_o_tag_ready[124]                  =   1'b0;
assign   tb_o_tag[124]                        =   tb_o_tag[123];

// CLK no. 125/1240
// *************************************************
assign   tb_i_valid[125]                      =   1'b0;
assign   tb_i_reset[125]                      =   1'b0;
assign   tb_i_sop[125]                        =   1'b0;
assign   tb_i_key_update[125]                 =   1'b0;
assign   tb_i_key[125]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[125]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[125]               =   1'b0;
assign   tb_i_rf_static_encrypt[125]          =   1'b1;
assign   tb_i_clear_fault_flags[125]          =   1'b0;
assign   tb_i_rf_static_aad_length[125]       =   64'h0000000000000100;
assign   tb_i_aad[125]                        =   tb_i_aad[124];
assign   tb_i_rf_static_plaintext_length[125] =   64'h0000000000000280;
assign   tb_i_plaintext[125]                  =   tb_i_plaintext[124];
assign   tb_o_valid[125]                      =   1'b0;
assign   tb_o_sop[125]                        =   1'b0;
assign   tb_o_ciphertext[125]                 =   tb_o_ciphertext[124];
assign   tb_o_tag_ready[125]                  =   1'b0;
assign   tb_o_tag[125]                        =   tb_o_tag[124];

// CLK no. 126/1240
// *************************************************
assign   tb_i_valid[126]                      =   1'b0;
assign   tb_i_reset[126]                      =   1'b0;
assign   tb_i_sop[126]                        =   1'b0;
assign   tb_i_key_update[126]                 =   1'b0;
assign   tb_i_key[126]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[126]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[126]               =   1'b0;
assign   tb_i_rf_static_encrypt[126]          =   1'b1;
assign   tb_i_clear_fault_flags[126]          =   1'b0;
assign   tb_i_rf_static_aad_length[126]       =   64'h0000000000000100;
assign   tb_i_aad[126]                        =   tb_i_aad[125];
assign   tb_i_rf_static_plaintext_length[126] =   64'h0000000000000280;
assign   tb_i_plaintext[126]                  =   tb_i_plaintext[125];
assign   tb_o_valid[126]                      =   1'b0;
assign   tb_o_sop[126]                        =   1'b0;
assign   tb_o_ciphertext[126]                 =   tb_o_ciphertext[125];
assign   tb_o_tag_ready[126]                  =   1'b0;
assign   tb_o_tag[126]                        =   tb_o_tag[125];

// CLK no. 127/1240
// *************************************************
assign   tb_i_valid[127]                      =   1'b0;
assign   tb_i_reset[127]                      =   1'b0;
assign   tb_i_sop[127]                        =   1'b0;
assign   tb_i_key_update[127]                 =   1'b0;
assign   tb_i_key[127]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[127]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[127]               =   1'b0;
assign   tb_i_rf_static_encrypt[127]          =   1'b1;
assign   tb_i_clear_fault_flags[127]          =   1'b0;
assign   tb_i_rf_static_aad_length[127]       =   64'h0000000000000100;
assign   tb_i_aad[127]                        =   tb_i_aad[126];
assign   tb_i_rf_static_plaintext_length[127] =   64'h0000000000000280;
assign   tb_i_plaintext[127]                  =   tb_i_plaintext[126];
assign   tb_o_valid[127]                      =   1'b0;
assign   tb_o_sop[127]                        =   1'b0;
assign   tb_o_ciphertext[127]                 =   tb_o_ciphertext[126];
assign   tb_o_tag_ready[127]                  =   1'b0;
assign   tb_o_tag[127]                        =   tb_o_tag[126];

// CLK no. 128/1240
// *************************************************
assign   tb_i_valid[128]                      =   1'b0;
assign   tb_i_reset[128]                      =   1'b0;
assign   tb_i_sop[128]                        =   1'b0;
assign   tb_i_key_update[128]                 =   1'b0;
assign   tb_i_key[128]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[128]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[128]               =   1'b0;
assign   tb_i_rf_static_encrypt[128]          =   1'b1;
assign   tb_i_clear_fault_flags[128]          =   1'b0;
assign   tb_i_rf_static_aad_length[128]       =   64'h0000000000000100;
assign   tb_i_aad[128]                        =   tb_i_aad[127];
assign   tb_i_rf_static_plaintext_length[128] =   64'h0000000000000280;
assign   tb_i_plaintext[128]                  =   tb_i_plaintext[127];
assign   tb_o_valid[128]                      =   1'b0;
assign   tb_o_sop[128]                        =   1'b0;
assign   tb_o_ciphertext[128]                 =   tb_o_ciphertext[127];
assign   tb_o_tag_ready[128]                  =   1'b0;
assign   tb_o_tag[128]                        =   tb_o_tag[127];

// CLK no. 129/1240
// *************************************************
assign   tb_i_valid[129]                      =   1'b0;
assign   tb_i_reset[129]                      =   1'b0;
assign   tb_i_sop[129]                        =   1'b0;
assign   tb_i_key_update[129]                 =   1'b0;
assign   tb_i_key[129]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[129]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[129]               =   1'b0;
assign   tb_i_rf_static_encrypt[129]          =   1'b1;
assign   tb_i_clear_fault_flags[129]          =   1'b0;
assign   tb_i_rf_static_aad_length[129]       =   64'h0000000000000100;
assign   tb_i_aad[129]                        =   tb_i_aad[128];
assign   tb_i_rf_static_plaintext_length[129] =   64'h0000000000000280;
assign   tb_i_plaintext[129]                  =   tb_i_plaintext[128];
assign   tb_o_valid[129]                      =   1'b0;
assign   tb_o_sop[129]                        =   1'b0;
assign   tb_o_ciphertext[129]                 =   tb_o_ciphertext[128];
assign   tb_o_tag_ready[129]                  =   1'b0;
assign   tb_o_tag[129]                        =   tb_o_tag[128];

// CLK no. 130/1240
// *************************************************
assign   tb_i_valid[130]                      =   1'b0;
assign   tb_i_reset[130]                      =   1'b0;
assign   tb_i_sop[130]                        =   1'b0;
assign   tb_i_key_update[130]                 =   1'b0;
assign   tb_i_key[130]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[130]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[130]               =   1'b0;
assign   tb_i_rf_static_encrypt[130]          =   1'b1;
assign   tb_i_clear_fault_flags[130]          =   1'b0;
assign   tb_i_rf_static_aad_length[130]       =   64'h0000000000000100;
assign   tb_i_aad[130]                        =   tb_i_aad[129];
assign   tb_i_rf_static_plaintext_length[130] =   64'h0000000000000280;
assign   tb_i_plaintext[130]                  =   tb_i_plaintext[129];
assign   tb_o_valid[130]                      =   1'b0;
assign   tb_o_sop[130]                        =   1'b0;
assign   tb_o_ciphertext[130]                 =   tb_o_ciphertext[129];
assign   tb_o_tag_ready[130]                  =   1'b0;
assign   tb_o_tag[130]                        =   tb_o_tag[129];

// CLK no. 131/1240
// *************************************************
assign   tb_i_valid[131]                      =   1'b0;
assign   tb_i_reset[131]                      =   1'b0;
assign   tb_i_sop[131]                        =   1'b0;
assign   tb_i_key_update[131]                 =   1'b0;
assign   tb_i_key[131]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[131]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[131]               =   1'b0;
assign   tb_i_rf_static_encrypt[131]          =   1'b1;
assign   tb_i_clear_fault_flags[131]          =   1'b0;
assign   tb_i_rf_static_aad_length[131]       =   64'h0000000000000100;
assign   tb_i_aad[131]                        =   tb_i_aad[130];
assign   tb_i_rf_static_plaintext_length[131] =   64'h0000000000000280;
assign   tb_i_plaintext[131]                  =   tb_i_plaintext[130];
assign   tb_o_valid[131]                      =   1'b0;
assign   tb_o_sop[131]                        =   1'b0;
assign   tb_o_ciphertext[131]                 =   tb_o_ciphertext[130];
assign   tb_o_tag_ready[131]                  =   1'b0;
assign   tb_o_tag[131]                        =   tb_o_tag[130];

// CLK no. 132/1240
// *************************************************
assign   tb_i_valid[132]                      =   1'b0;
assign   tb_i_reset[132]                      =   1'b0;
assign   tb_i_sop[132]                        =   1'b0;
assign   tb_i_key_update[132]                 =   1'b0;
assign   tb_i_key[132]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[132]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[132]               =   1'b0;
assign   tb_i_rf_static_encrypt[132]          =   1'b1;
assign   tb_i_clear_fault_flags[132]          =   1'b0;
assign   tb_i_rf_static_aad_length[132]       =   64'h0000000000000100;
assign   tb_i_aad[132]                        =   tb_i_aad[131];
assign   tb_i_rf_static_plaintext_length[132] =   64'h0000000000000280;
assign   tb_i_plaintext[132]                  =   tb_i_plaintext[131];
assign   tb_o_valid[132]                      =   1'b0;
assign   tb_o_sop[132]                        =   1'b0;
assign   tb_o_ciphertext[132]                 =   tb_o_ciphertext[131];
assign   tb_o_tag_ready[132]                  =   1'b0;
assign   tb_o_tag[132]                        =   tb_o_tag[131];

// CLK no. 133/1240
// *************************************************
assign   tb_i_valid[133]                      =   1'b0;
assign   tb_i_reset[133]                      =   1'b0;
assign   tb_i_sop[133]                        =   1'b0;
assign   tb_i_key_update[133]                 =   1'b0;
assign   tb_i_key[133]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[133]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[133]               =   1'b0;
assign   tb_i_rf_static_encrypt[133]          =   1'b1;
assign   tb_i_clear_fault_flags[133]          =   1'b0;
assign   tb_i_rf_static_aad_length[133]       =   64'h0000000000000100;
assign   tb_i_aad[133]                        =   tb_i_aad[132];
assign   tb_i_rf_static_plaintext_length[133] =   64'h0000000000000280;
assign   tb_i_plaintext[133]                  =   tb_i_plaintext[132];
assign   tb_o_valid[133]                      =   1'b0;
assign   tb_o_sop[133]                        =   1'b0;
assign   tb_o_ciphertext[133]                 =   tb_o_ciphertext[132];
assign   tb_o_tag_ready[133]                  =   1'b0;
assign   tb_o_tag[133]                        =   tb_o_tag[132];

// CLK no. 134/1240
// *************************************************
assign   tb_i_valid[134]                      =   1'b0;
assign   tb_i_reset[134]                      =   1'b0;
assign   tb_i_sop[134]                        =   1'b0;
assign   tb_i_key_update[134]                 =   1'b0;
assign   tb_i_key[134]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[134]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[134]               =   1'b0;
assign   tb_i_rf_static_encrypt[134]          =   1'b1;
assign   tb_i_clear_fault_flags[134]          =   1'b0;
assign   tb_i_rf_static_aad_length[134]       =   64'h0000000000000100;
assign   tb_i_aad[134]                        =   tb_i_aad[133];
assign   tb_i_rf_static_plaintext_length[134] =   64'h0000000000000280;
assign   tb_i_plaintext[134]                  =   tb_i_plaintext[133];
assign   tb_o_valid[134]                      =   1'b0;
assign   tb_o_sop[134]                        =   1'b0;
assign   tb_o_ciphertext[134]                 =   tb_o_ciphertext[133];
assign   tb_o_tag_ready[134]                  =   1'b0;
assign   tb_o_tag[134]                        =   tb_o_tag[133];

// CLK no. 135/1240
// *************************************************
assign   tb_i_valid[135]                      =   1'b0;
assign   tb_i_reset[135]                      =   1'b0;
assign   tb_i_sop[135]                        =   1'b0;
assign   tb_i_key_update[135]                 =   1'b0;
assign   tb_i_key[135]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[135]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[135]               =   1'b0;
assign   tb_i_rf_static_encrypt[135]          =   1'b1;
assign   tb_i_clear_fault_flags[135]          =   1'b0;
assign   tb_i_rf_static_aad_length[135]       =   64'h0000000000000100;
assign   tb_i_aad[135]                        =   tb_i_aad[134];
assign   tb_i_rf_static_plaintext_length[135] =   64'h0000000000000280;
assign   tb_i_plaintext[135]                  =   tb_i_plaintext[134];
assign   tb_o_valid[135]                      =   1'b0;
assign   tb_o_sop[135]                        =   1'b0;
assign   tb_o_ciphertext[135]                 =   tb_o_ciphertext[134];
assign   tb_o_tag_ready[135]                  =   1'b0;
assign   tb_o_tag[135]                        =   tb_o_tag[134];

// CLK no. 136/1240
// *************************************************
assign   tb_i_valid[136]                      =   1'b0;
assign   tb_i_reset[136]                      =   1'b0;
assign   tb_i_sop[136]                        =   1'b0;
assign   tb_i_key_update[136]                 =   1'b0;
assign   tb_i_key[136]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[136]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[136]               =   1'b0;
assign   tb_i_rf_static_encrypt[136]          =   1'b1;
assign   tb_i_clear_fault_flags[136]          =   1'b0;
assign   tb_i_rf_static_aad_length[136]       =   64'h0000000000000100;
assign   tb_i_aad[136]                        =   tb_i_aad[135];
assign   tb_i_rf_static_plaintext_length[136] =   64'h0000000000000280;
assign   tb_i_plaintext[136]                  =   tb_i_plaintext[135];
assign   tb_o_valid[136]                      =   1'b0;
assign   tb_o_sop[136]                        =   1'b0;
assign   tb_o_ciphertext[136]                 =   tb_o_ciphertext[135];
assign   tb_o_tag_ready[136]                  =   1'b0;
assign   tb_o_tag[136]                        =   tb_o_tag[135];

// CLK no. 137/1240
// *************************************************
assign   tb_i_valid[137]                      =   1'b0;
assign   tb_i_reset[137]                      =   1'b0;
assign   tb_i_sop[137]                        =   1'b0;
assign   tb_i_key_update[137]                 =   1'b0;
assign   tb_i_key[137]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[137]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[137]               =   1'b0;
assign   tb_i_rf_static_encrypt[137]          =   1'b1;
assign   tb_i_clear_fault_flags[137]          =   1'b0;
assign   tb_i_rf_static_aad_length[137]       =   64'h0000000000000100;
assign   tb_i_aad[137]                        =   tb_i_aad[136];
assign   tb_i_rf_static_plaintext_length[137] =   64'h0000000000000280;
assign   tb_i_plaintext[137]                  =   tb_i_plaintext[136];
assign   tb_o_valid[137]                      =   1'b0;
assign   tb_o_sop[137]                        =   1'b0;
assign   tb_o_ciphertext[137]                 =   tb_o_ciphertext[136];
assign   tb_o_tag_ready[137]                  =   1'b0;
assign   tb_o_tag[137]                        =   tb_o_tag[136];

// CLK no. 138/1240
// *************************************************
assign   tb_i_valid[138]                      =   1'b0;
assign   tb_i_reset[138]                      =   1'b0;
assign   tb_i_sop[138]                        =   1'b0;
assign   tb_i_key_update[138]                 =   1'b0;
assign   tb_i_key[138]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[138]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[138]               =   1'b0;
assign   tb_i_rf_static_encrypt[138]          =   1'b1;
assign   tb_i_clear_fault_flags[138]          =   1'b0;
assign   tb_i_rf_static_aad_length[138]       =   64'h0000000000000100;
assign   tb_i_aad[138]                        =   tb_i_aad[137];
assign   tb_i_rf_static_plaintext_length[138] =   64'h0000000000000280;
assign   tb_i_plaintext[138]                  =   tb_i_plaintext[137];
assign   tb_o_valid[138]                      =   1'b0;
assign   tb_o_sop[138]                        =   1'b0;
assign   tb_o_ciphertext[138]                 =   tb_o_ciphertext[137];
assign   tb_o_tag_ready[138]                  =   1'b0;
assign   tb_o_tag[138]                        =   tb_o_tag[137];

// CLK no. 139/1240
// *************************************************
assign   tb_i_valid[139]                      =   1'b0;
assign   tb_i_reset[139]                      =   1'b0;
assign   tb_i_sop[139]                        =   1'b0;
assign   tb_i_key_update[139]                 =   1'b0;
assign   tb_i_key[139]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[139]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[139]               =   1'b0;
assign   tb_i_rf_static_encrypt[139]          =   1'b1;
assign   tb_i_clear_fault_flags[139]          =   1'b0;
assign   tb_i_rf_static_aad_length[139]       =   64'h0000000000000100;
assign   tb_i_aad[139]                        =   tb_i_aad[138];
assign   tb_i_rf_static_plaintext_length[139] =   64'h0000000000000280;
assign   tb_i_plaintext[139]                  =   tb_i_plaintext[138];
assign   tb_o_valid[139]                      =   1'b0;
assign   tb_o_sop[139]                        =   1'b0;
assign   tb_o_ciphertext[139]                 =   tb_o_ciphertext[138];
assign   tb_o_tag_ready[139]                  =   1'b0;
assign   tb_o_tag[139]                        =   tb_o_tag[138];

// CLK no. 140/1240
// *************************************************
assign   tb_i_valid[140]                      =   1'b0;
assign   tb_i_reset[140]                      =   1'b0;
assign   tb_i_sop[140]                        =   1'b0;
assign   tb_i_key_update[140]                 =   1'b0;
assign   tb_i_key[140]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[140]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[140]               =   1'b0;
assign   tb_i_rf_static_encrypt[140]          =   1'b1;
assign   tb_i_clear_fault_flags[140]          =   1'b0;
assign   tb_i_rf_static_aad_length[140]       =   64'h0000000000000100;
assign   tb_i_aad[140]                        =   tb_i_aad[139];
assign   tb_i_rf_static_plaintext_length[140] =   64'h0000000000000280;
assign   tb_i_plaintext[140]                  =   tb_i_plaintext[139];
assign   tb_o_valid[140]                      =   1'b0;
assign   tb_o_sop[140]                        =   1'b0;
assign   tb_o_ciphertext[140]                 =   tb_o_ciphertext[139];
assign   tb_o_tag_ready[140]                  =   1'b0;
assign   tb_o_tag[140]                        =   tb_o_tag[139];

// CLK no. 141/1240
// *************************************************
assign   tb_i_valid[141]                      =   1'b0;
assign   tb_i_reset[141]                      =   1'b0;
assign   tb_i_sop[141]                        =   1'b0;
assign   tb_i_key_update[141]                 =   1'b0;
assign   tb_i_key[141]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[141]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[141]               =   1'b0;
assign   tb_i_rf_static_encrypt[141]          =   1'b1;
assign   tb_i_clear_fault_flags[141]          =   1'b0;
assign   tb_i_rf_static_aad_length[141]       =   64'h0000000000000100;
assign   tb_i_aad[141]                        =   tb_i_aad[140];
assign   tb_i_rf_static_plaintext_length[141] =   64'h0000000000000280;
assign   tb_i_plaintext[141]                  =   tb_i_plaintext[140];
assign   tb_o_valid[141]                      =   1'b0;
assign   tb_o_sop[141]                        =   1'b0;
assign   tb_o_ciphertext[141]                 =   tb_o_ciphertext[140];
assign   tb_o_tag_ready[141]                  =   1'b0;
assign   tb_o_tag[141]                        =   tb_o_tag[140];

// CLK no. 142/1240
// *************************************************
assign   tb_i_valid[142]                      =   1'b0;
assign   tb_i_reset[142]                      =   1'b0;
assign   tb_i_sop[142]                        =   1'b0;
assign   tb_i_key_update[142]                 =   1'b0;
assign   tb_i_key[142]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[142]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[142]               =   1'b0;
assign   tb_i_rf_static_encrypt[142]          =   1'b1;
assign   tb_i_clear_fault_flags[142]          =   1'b0;
assign   tb_i_rf_static_aad_length[142]       =   64'h0000000000000100;
assign   tb_i_aad[142]                        =   tb_i_aad[141];
assign   tb_i_rf_static_plaintext_length[142] =   64'h0000000000000280;
assign   tb_i_plaintext[142]                  =   tb_i_plaintext[141];
assign   tb_o_valid[142]                      =   1'b0;
assign   tb_o_sop[142]                        =   1'b0;
assign   tb_o_ciphertext[142]                 =   tb_o_ciphertext[141];
assign   tb_o_tag_ready[142]                  =   1'b0;
assign   tb_o_tag[142]                        =   tb_o_tag[141];

// CLK no. 143/1240
// *************************************************
assign   tb_i_valid[143]                      =   1'b0;
assign   tb_i_reset[143]                      =   1'b0;
assign   tb_i_sop[143]                        =   1'b0;
assign   tb_i_key_update[143]                 =   1'b0;
assign   tb_i_key[143]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[143]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[143]               =   1'b0;
assign   tb_i_rf_static_encrypt[143]          =   1'b1;
assign   tb_i_clear_fault_flags[143]          =   1'b0;
assign   tb_i_rf_static_aad_length[143]       =   64'h0000000000000100;
assign   tb_i_aad[143]                        =   tb_i_aad[142];
assign   tb_i_rf_static_plaintext_length[143] =   64'h0000000000000280;
assign   tb_i_plaintext[143]                  =   tb_i_plaintext[142];
assign   tb_o_valid[143]                      =   1'b0;
assign   tb_o_sop[143]                        =   1'b0;
assign   tb_o_ciphertext[143]                 =   tb_o_ciphertext[142];
assign   tb_o_tag_ready[143]                  =   1'b0;
assign   tb_o_tag[143]                        =   tb_o_tag[142];

// CLK no. 144/1240
// *************************************************
assign   tb_i_valid[144]                      =   1'b0;
assign   tb_i_reset[144]                      =   1'b0;
assign   tb_i_sop[144]                        =   1'b0;
assign   tb_i_key_update[144]                 =   1'b0;
assign   tb_i_key[144]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[144]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[144]               =   1'b0;
assign   tb_i_rf_static_encrypt[144]          =   1'b1;
assign   tb_i_clear_fault_flags[144]          =   1'b0;
assign   tb_i_rf_static_aad_length[144]       =   64'h0000000000000100;
assign   tb_i_aad[144]                        =   tb_i_aad[143];
assign   tb_i_rf_static_plaintext_length[144] =   64'h0000000000000280;
assign   tb_i_plaintext[144]                  =   tb_i_plaintext[143];
assign   tb_o_valid[144]                      =   1'b0;
assign   tb_o_sop[144]                        =   1'b0;
assign   tb_o_ciphertext[144]                 =   tb_o_ciphertext[143];
assign   tb_o_tag_ready[144]                  =   1'b0;
assign   tb_o_tag[144]                        =   tb_o_tag[143];

// CLK no. 145/1240
// *************************************************
assign   tb_i_valid[145]                      =   1'b0;
assign   tb_i_reset[145]                      =   1'b0;
assign   tb_i_sop[145]                        =   1'b0;
assign   tb_i_key_update[145]                 =   1'b0;
assign   tb_i_key[145]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[145]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[145]               =   1'b0;
assign   tb_i_rf_static_encrypt[145]          =   1'b1;
assign   tb_i_clear_fault_flags[145]          =   1'b0;
assign   tb_i_rf_static_aad_length[145]       =   64'h0000000000000100;
assign   tb_i_aad[145]                        =   tb_i_aad[144];
assign   tb_i_rf_static_plaintext_length[145] =   64'h0000000000000280;
assign   tb_i_plaintext[145]                  =   tb_i_plaintext[144];
assign   tb_o_valid[145]                      =   1'b0;
assign   tb_o_sop[145]                        =   1'b0;
assign   tb_o_ciphertext[145]                 =   tb_o_ciphertext[144];
assign   tb_o_tag_ready[145]                  =   1'b0;
assign   tb_o_tag[145]                        =   tb_o_tag[144];

// CLK no. 146/1240
// *************************************************
assign   tb_i_valid[146]                      =   1'b0;
assign   tb_i_reset[146]                      =   1'b0;
assign   tb_i_sop[146]                        =   1'b0;
assign   tb_i_key_update[146]                 =   1'b0;
assign   tb_i_key[146]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[146]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[146]               =   1'b0;
assign   tb_i_rf_static_encrypt[146]          =   1'b1;
assign   tb_i_clear_fault_flags[146]          =   1'b0;
assign   tb_i_rf_static_aad_length[146]       =   64'h0000000000000100;
assign   tb_i_aad[146]                        =   tb_i_aad[145];
assign   tb_i_rf_static_plaintext_length[146] =   64'h0000000000000280;
assign   tb_i_plaintext[146]                  =   tb_i_plaintext[145];
assign   tb_o_valid[146]                      =   1'b0;
assign   tb_o_sop[146]                        =   1'b0;
assign   tb_o_ciphertext[146]                 =   tb_o_ciphertext[145];
assign   tb_o_tag_ready[146]                  =   1'b0;
assign   tb_o_tag[146]                        =   tb_o_tag[145];

// CLK no. 147/1240
// *************************************************
assign   tb_i_valid[147]                      =   1'b0;
assign   tb_i_reset[147]                      =   1'b0;
assign   tb_i_sop[147]                        =   1'b0;
assign   tb_i_key_update[147]                 =   1'b0;
assign   tb_i_key[147]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[147]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[147]               =   1'b0;
assign   tb_i_rf_static_encrypt[147]          =   1'b1;
assign   tb_i_clear_fault_flags[147]          =   1'b0;
assign   tb_i_rf_static_aad_length[147]       =   64'h0000000000000100;
assign   tb_i_aad[147]                        =   tb_i_aad[146];
assign   tb_i_rf_static_plaintext_length[147] =   64'h0000000000000280;
assign   tb_i_plaintext[147]                  =   tb_i_plaintext[146];
assign   tb_o_valid[147]                      =   1'b0;
assign   tb_o_sop[147]                        =   1'b0;
assign   tb_o_ciphertext[147]                 =   tb_o_ciphertext[146];
assign   tb_o_tag_ready[147]                  =   1'b0;
assign   tb_o_tag[147]                        =   tb_o_tag[146];

// CLK no. 148/1240
// *************************************************
assign   tb_i_valid[148]                      =   1'b0;
assign   tb_i_reset[148]                      =   1'b0;
assign   tb_i_sop[148]                        =   1'b0;
assign   tb_i_key_update[148]                 =   1'b0;
assign   tb_i_key[148]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[148]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[148]               =   1'b0;
assign   tb_i_rf_static_encrypt[148]          =   1'b1;
assign   tb_i_clear_fault_flags[148]          =   1'b0;
assign   tb_i_rf_static_aad_length[148]       =   64'h0000000000000100;
assign   tb_i_aad[148]                        =   tb_i_aad[147];
assign   tb_i_rf_static_plaintext_length[148] =   64'h0000000000000280;
assign   tb_i_plaintext[148]                  =   tb_i_plaintext[147];
assign   tb_o_valid[148]                      =   1'b0;
assign   tb_o_sop[148]                        =   1'b0;
assign   tb_o_ciphertext[148]                 =   tb_o_ciphertext[147];
assign   tb_o_tag_ready[148]                  =   1'b0;
assign   tb_o_tag[148]                        =   tb_o_tag[147];

// CLK no. 149/1240
// *************************************************
assign   tb_i_valid[149]                      =   1'b0;
assign   tb_i_reset[149]                      =   1'b0;
assign   tb_i_sop[149]                        =   1'b0;
assign   tb_i_key_update[149]                 =   1'b0;
assign   tb_i_key[149]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[149]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[149]               =   1'b0;
assign   tb_i_rf_static_encrypt[149]          =   1'b1;
assign   tb_i_clear_fault_flags[149]          =   1'b0;
assign   tb_i_rf_static_aad_length[149]       =   64'h0000000000000100;
assign   tb_i_aad[149]                        =   tb_i_aad[148];
assign   tb_i_rf_static_plaintext_length[149] =   64'h0000000000000280;
assign   tb_i_plaintext[149]                  =   tb_i_plaintext[148];
assign   tb_o_valid[149]                      =   1'b0;
assign   tb_o_sop[149]                        =   1'b0;
assign   tb_o_ciphertext[149]                 =   tb_o_ciphertext[148];
assign   tb_o_tag_ready[149]                  =   1'b0;
assign   tb_o_tag[149]                        =   tb_o_tag[148];

// CLK no. 150/1240
// *************************************************
assign   tb_i_valid[150]                      =   1'b0;
assign   tb_i_reset[150]                      =   1'b0;
assign   tb_i_sop[150]                        =   1'b0;
assign   tb_i_key_update[150]                 =   1'b0;
assign   tb_i_key[150]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[150]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[150]               =   1'b0;
assign   tb_i_rf_static_encrypt[150]          =   1'b1;
assign   tb_i_clear_fault_flags[150]          =   1'b0;
assign   tb_i_rf_static_aad_length[150]       =   64'h0000000000000100;
assign   tb_i_aad[150]                        =   tb_i_aad[149];
assign   tb_i_rf_static_plaintext_length[150] =   64'h0000000000000280;
assign   tb_i_plaintext[150]                  =   tb_i_plaintext[149];
assign   tb_o_valid[150]                      =   1'b0;
assign   tb_o_sop[150]                        =   1'b0;
assign   tb_o_ciphertext[150]                 =   tb_o_ciphertext[149];
assign   tb_o_tag_ready[150]                  =   1'b0;
assign   tb_o_tag[150]                        =   tb_o_tag[149];

// CLK no. 151/1240
// *************************************************
assign   tb_i_valid[151]                      =   1'b0;
assign   tb_i_reset[151]                      =   1'b0;
assign   tb_i_sop[151]                        =   1'b0;
assign   tb_i_key_update[151]                 =   1'b0;
assign   tb_i_key[151]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[151]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[151]               =   1'b0;
assign   tb_i_rf_static_encrypt[151]          =   1'b1;
assign   tb_i_clear_fault_flags[151]          =   1'b0;
assign   tb_i_rf_static_aad_length[151]       =   64'h0000000000000100;
assign   tb_i_aad[151]                        =   tb_i_aad[150];
assign   tb_i_rf_static_plaintext_length[151] =   64'h0000000000000280;
assign   tb_i_plaintext[151]                  =   tb_i_plaintext[150];
assign   tb_o_valid[151]                      =   1'b0;
assign   tb_o_sop[151]                        =   1'b0;
assign   tb_o_ciphertext[151]                 =   tb_o_ciphertext[150];
assign   tb_o_tag_ready[151]                  =   1'b0;
assign   tb_o_tag[151]                        =   tb_o_tag[150];

// CLK no. 152/1240
// *************************************************
assign   tb_i_valid[152]                      =   1'b0;
assign   tb_i_reset[152]                      =   1'b0;
assign   tb_i_sop[152]                        =   1'b0;
assign   tb_i_key_update[152]                 =   1'b0;
assign   tb_i_key[152]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[152]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[152]               =   1'b0;
assign   tb_i_rf_static_encrypt[152]          =   1'b1;
assign   tb_i_clear_fault_flags[152]          =   1'b0;
assign   tb_i_rf_static_aad_length[152]       =   64'h0000000000000100;
assign   tb_i_aad[152]                        =   tb_i_aad[151];
assign   tb_i_rf_static_plaintext_length[152] =   64'h0000000000000280;
assign   tb_i_plaintext[152]                  =   tb_i_plaintext[151];
assign   tb_o_valid[152]                      =   1'b0;
assign   tb_o_sop[152]                        =   1'b0;
assign   tb_o_ciphertext[152]                 =   tb_o_ciphertext[151];
assign   tb_o_tag_ready[152]                  =   1'b0;
assign   tb_o_tag[152]                        =   tb_o_tag[151];

// CLK no. 153/1240
// *************************************************
assign   tb_i_valid[153]                      =   1'b0;
assign   tb_i_reset[153]                      =   1'b0;
assign   tb_i_sop[153]                        =   1'b0;
assign   tb_i_key_update[153]                 =   1'b0;
assign   tb_i_key[153]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[153]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[153]               =   1'b0;
assign   tb_i_rf_static_encrypt[153]          =   1'b1;
assign   tb_i_clear_fault_flags[153]          =   1'b0;
assign   tb_i_rf_static_aad_length[153]       =   64'h0000000000000100;
assign   tb_i_aad[153]                        =   tb_i_aad[152];
assign   tb_i_rf_static_plaintext_length[153] =   64'h0000000000000280;
assign   tb_i_plaintext[153]                  =   tb_i_plaintext[152];
assign   tb_o_valid[153]                      =   1'b0;
assign   tb_o_sop[153]                        =   1'b0;
assign   tb_o_ciphertext[153]                 =   tb_o_ciphertext[152];
assign   tb_o_tag_ready[153]                  =   1'b0;
assign   tb_o_tag[153]                        =   tb_o_tag[152];

// CLK no. 154/1240
// *************************************************
assign   tb_i_valid[154]                      =   1'b0;
assign   tb_i_reset[154]                      =   1'b0;
assign   tb_i_sop[154]                        =   1'b0;
assign   tb_i_key_update[154]                 =   1'b0;
assign   tb_i_key[154]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[154]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[154]               =   1'b0;
assign   tb_i_rf_static_encrypt[154]          =   1'b1;
assign   tb_i_clear_fault_flags[154]          =   1'b0;
assign   tb_i_rf_static_aad_length[154]       =   64'h0000000000000100;
assign   tb_i_aad[154]                        =   tb_i_aad[153];
assign   tb_i_rf_static_plaintext_length[154] =   64'h0000000000000280;
assign   tb_i_plaintext[154]                  =   tb_i_plaintext[153];
assign   tb_o_valid[154]                      =   1'b0;
assign   tb_o_sop[154]                        =   1'b0;
assign   tb_o_ciphertext[154]                 =   tb_o_ciphertext[153];
assign   tb_o_tag_ready[154]                  =   1'b0;
assign   tb_o_tag[154]                        =   tb_o_tag[153];

// CLK no. 155/1240
// *************************************************
assign   tb_i_valid[155]                      =   1'b0;
assign   tb_i_reset[155]                      =   1'b0;
assign   tb_i_sop[155]                        =   1'b0;
assign   tb_i_key_update[155]                 =   1'b0;
assign   tb_i_key[155]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[155]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[155]               =   1'b0;
assign   tb_i_rf_static_encrypt[155]          =   1'b1;
assign   tb_i_clear_fault_flags[155]          =   1'b0;
assign   tb_i_rf_static_aad_length[155]       =   64'h0000000000000100;
assign   tb_i_aad[155]                        =   tb_i_aad[154];
assign   tb_i_rf_static_plaintext_length[155] =   64'h0000000000000280;
assign   tb_i_plaintext[155]                  =   tb_i_plaintext[154];
assign   tb_o_valid[155]                      =   1'b0;
assign   tb_o_sop[155]                        =   1'b0;
assign   tb_o_ciphertext[155]                 =   tb_o_ciphertext[154];
assign   tb_o_tag_ready[155]                  =   1'b0;
assign   tb_o_tag[155]                        =   tb_o_tag[154];

// CLK no. 156/1240
// *************************************************
assign   tb_i_valid[156]                      =   1'b0;
assign   tb_i_reset[156]                      =   1'b0;
assign   tb_i_sop[156]                        =   1'b0;
assign   tb_i_key_update[156]                 =   1'b0;
assign   tb_i_key[156]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[156]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[156]               =   1'b0;
assign   tb_i_rf_static_encrypt[156]          =   1'b1;
assign   tb_i_clear_fault_flags[156]          =   1'b0;
assign   tb_i_rf_static_aad_length[156]       =   64'h0000000000000100;
assign   tb_i_aad[156]                        =   tb_i_aad[155];
assign   tb_i_rf_static_plaintext_length[156] =   64'h0000000000000280;
assign   tb_i_plaintext[156]                  =   tb_i_plaintext[155];
assign   tb_o_valid[156]                      =   1'b0;
assign   tb_o_sop[156]                        =   1'b0;
assign   tb_o_ciphertext[156]                 =   tb_o_ciphertext[155];
assign   tb_o_tag_ready[156]                  =   1'b0;
assign   tb_o_tag[156]                        =   tb_o_tag[155];

// CLK no. 157/1240
// *************************************************
assign   tb_i_valid[157]                      =   1'b0;
assign   tb_i_reset[157]                      =   1'b0;
assign   tb_i_sop[157]                        =   1'b0;
assign   tb_i_key_update[157]                 =   1'b0;
assign   tb_i_key[157]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[157]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[157]               =   1'b0;
assign   tb_i_rf_static_encrypt[157]          =   1'b1;
assign   tb_i_clear_fault_flags[157]          =   1'b0;
assign   tb_i_rf_static_aad_length[157]       =   64'h0000000000000100;
assign   tb_i_aad[157]                        =   tb_i_aad[156];
assign   tb_i_rf_static_plaintext_length[157] =   64'h0000000000000280;
assign   tb_i_plaintext[157]                  =   tb_i_plaintext[156];
assign   tb_o_valid[157]                      =   1'b0;
assign   tb_o_sop[157]                        =   1'b0;
assign   tb_o_ciphertext[157]                 =   tb_o_ciphertext[156];
assign   tb_o_tag_ready[157]                  =   1'b0;
assign   tb_o_tag[157]                        =   tb_o_tag[156];

// CLK no. 158/1240
// *************************************************
assign   tb_i_valid[158]                      =   1'b0;
assign   tb_i_reset[158]                      =   1'b0;
assign   tb_i_sop[158]                        =   1'b0;
assign   tb_i_key_update[158]                 =   1'b0;
assign   tb_i_key[158]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[158]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[158]               =   1'b0;
assign   tb_i_rf_static_encrypt[158]          =   1'b1;
assign   tb_i_clear_fault_flags[158]          =   1'b0;
assign   tb_i_rf_static_aad_length[158]       =   64'h0000000000000100;
assign   tb_i_aad[158]                        =   tb_i_aad[157];
assign   tb_i_rf_static_plaintext_length[158] =   64'h0000000000000280;
assign   tb_i_plaintext[158]                  =   tb_i_plaintext[157];
assign   tb_o_valid[158]                      =   1'b0;
assign   tb_o_sop[158]                        =   1'b0;
assign   tb_o_ciphertext[158]                 =   tb_o_ciphertext[157];
assign   tb_o_tag_ready[158]                  =   1'b0;
assign   tb_o_tag[158]                        =   tb_o_tag[157];

// CLK no. 159/1240
// *************************************************
assign   tb_i_valid[159]                      =   1'b0;
assign   tb_i_reset[159]                      =   1'b0;
assign   tb_i_sop[159]                        =   1'b0;
assign   tb_i_key_update[159]                 =   1'b0;
assign   tb_i_key[159]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[159]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[159]               =   1'b0;
assign   tb_i_rf_static_encrypt[159]          =   1'b1;
assign   tb_i_clear_fault_flags[159]          =   1'b0;
assign   tb_i_rf_static_aad_length[159]       =   64'h0000000000000100;
assign   tb_i_aad[159]                        =   tb_i_aad[158];
assign   tb_i_rf_static_plaintext_length[159] =   64'h0000000000000280;
assign   tb_i_plaintext[159]                  =   tb_i_plaintext[158];
assign   tb_o_valid[159]                      =   1'b0;
assign   tb_o_sop[159]                        =   1'b0;
assign   tb_o_ciphertext[159]                 =   tb_o_ciphertext[158];
assign   tb_o_tag_ready[159]                  =   1'b0;
assign   tb_o_tag[159]                        =   tb_o_tag[158];

// CLK no. 160/1240
// *************************************************
assign   tb_i_valid[160]                      =   1'b0;
assign   tb_i_reset[160]                      =   1'b0;
assign   tb_i_sop[160]                        =   1'b0;
assign   tb_i_key_update[160]                 =   1'b0;
assign   tb_i_key[160]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[160]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[160]               =   1'b0;
assign   tb_i_rf_static_encrypt[160]          =   1'b1;
assign   tb_i_clear_fault_flags[160]          =   1'b0;
assign   tb_i_rf_static_aad_length[160]       =   64'h0000000000000100;
assign   tb_i_aad[160]                        =   tb_i_aad[159];
assign   tb_i_rf_static_plaintext_length[160] =   64'h0000000000000280;
assign   tb_i_plaintext[160]                  =   tb_i_plaintext[159];
assign   tb_o_valid[160]                      =   1'b0;
assign   tb_o_sop[160]                        =   1'b0;
assign   tb_o_ciphertext[160]                 =   tb_o_ciphertext[159];
assign   tb_o_tag_ready[160]                  =   1'b0;
assign   tb_o_tag[160]                        =   tb_o_tag[159];

// CLK no. 161/1240
// *************************************************
assign   tb_i_valid[161]                      =   1'b0;
assign   tb_i_reset[161]                      =   1'b0;
assign   tb_i_sop[161]                        =   1'b0;
assign   tb_i_key_update[161]                 =   1'b0;
assign   tb_i_key[161]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[161]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[161]               =   1'b0;
assign   tb_i_rf_static_encrypt[161]          =   1'b1;
assign   tb_i_clear_fault_flags[161]          =   1'b0;
assign   tb_i_rf_static_aad_length[161]       =   64'h0000000000000100;
assign   tb_i_aad[161]                        =   tb_i_aad[160];
assign   tb_i_rf_static_plaintext_length[161] =   64'h0000000000000280;
assign   tb_i_plaintext[161]                  =   tb_i_plaintext[160];
assign   tb_o_valid[161]                      =   1'b0;
assign   tb_o_sop[161]                        =   1'b0;
assign   tb_o_ciphertext[161]                 =   tb_o_ciphertext[160];
assign   tb_o_tag_ready[161]                  =   1'b0;
assign   tb_o_tag[161]                        =   tb_o_tag[160];

// CLK no. 162/1240
// *************************************************
assign   tb_i_valid[162]                      =   1'b0;
assign   tb_i_reset[162]                      =   1'b0;
assign   tb_i_sop[162]                        =   1'b0;
assign   tb_i_key_update[162]                 =   1'b0;
assign   tb_i_key[162]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[162]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[162]               =   1'b0;
assign   tb_i_rf_static_encrypt[162]          =   1'b1;
assign   tb_i_clear_fault_flags[162]          =   1'b0;
assign   tb_i_rf_static_aad_length[162]       =   64'h0000000000000100;
assign   tb_i_aad[162]                        =   tb_i_aad[161];
assign   tb_i_rf_static_plaintext_length[162] =   64'h0000000000000280;
assign   tb_i_plaintext[162]                  =   tb_i_plaintext[161];
assign   tb_o_valid[162]                      =   1'b0;
assign   tb_o_sop[162]                        =   1'b0;
assign   tb_o_ciphertext[162]                 =   tb_o_ciphertext[161];
assign   tb_o_tag_ready[162]                  =   1'b0;
assign   tb_o_tag[162]                        =   tb_o_tag[161];

// CLK no. 163/1240
// *************************************************
assign   tb_i_valid[163]                      =   1'b0;
assign   tb_i_reset[163]                      =   1'b0;
assign   tb_i_sop[163]                        =   1'b0;
assign   tb_i_key_update[163]                 =   1'b0;
assign   tb_i_key[163]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[163]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[163]               =   1'b0;
assign   tb_i_rf_static_encrypt[163]          =   1'b1;
assign   tb_i_clear_fault_flags[163]          =   1'b0;
assign   tb_i_rf_static_aad_length[163]       =   64'h0000000000000100;
assign   tb_i_aad[163]                        =   tb_i_aad[162];
assign   tb_i_rf_static_plaintext_length[163] =   64'h0000000000000280;
assign   tb_i_plaintext[163]                  =   tb_i_plaintext[162];
assign   tb_o_valid[163]                      =   1'b0;
assign   tb_o_sop[163]                        =   1'b0;
assign   tb_o_ciphertext[163]                 =   tb_o_ciphertext[162];
assign   tb_o_tag_ready[163]                  =   1'b0;
assign   tb_o_tag[163]                        =   tb_o_tag[162];

// CLK no. 164/1240
// *************************************************
assign   tb_i_valid[164]                      =   1'b0;
assign   tb_i_reset[164]                      =   1'b0;
assign   tb_i_sop[164]                        =   1'b0;
assign   tb_i_key_update[164]                 =   1'b0;
assign   tb_i_key[164]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[164]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[164]               =   1'b0;
assign   tb_i_rf_static_encrypt[164]          =   1'b1;
assign   tb_i_clear_fault_flags[164]          =   1'b0;
assign   tb_i_rf_static_aad_length[164]       =   64'h0000000000000100;
assign   tb_i_aad[164]                        =   tb_i_aad[163];
assign   tb_i_rf_static_plaintext_length[164] =   64'h0000000000000280;
assign   tb_i_plaintext[164]                  =   tb_i_plaintext[163];
assign   tb_o_valid[164]                      =   1'b0;
assign   tb_o_sop[164]                        =   1'b0;
assign   tb_o_ciphertext[164]                 =   tb_o_ciphertext[163];
assign   tb_o_tag_ready[164]                  =   1'b0;
assign   tb_o_tag[164]                        =   tb_o_tag[163];

// CLK no. 165/1240
// *************************************************
assign   tb_i_valid[165]                      =   1'b0;
assign   tb_i_reset[165]                      =   1'b0;
assign   tb_i_sop[165]                        =   1'b0;
assign   tb_i_key_update[165]                 =   1'b0;
assign   tb_i_key[165]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[165]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[165]               =   1'b0;
assign   tb_i_rf_static_encrypt[165]          =   1'b1;
assign   tb_i_clear_fault_flags[165]          =   1'b0;
assign   tb_i_rf_static_aad_length[165]       =   64'h0000000000000100;
assign   tb_i_aad[165]                        =   tb_i_aad[164];
assign   tb_i_rf_static_plaintext_length[165] =   64'h0000000000000280;
assign   tb_i_plaintext[165]                  =   tb_i_plaintext[164];
assign   tb_o_valid[165]                      =   1'b1;
assign   tb_o_sop[165]                        =   1'b1;
assign   tb_o_ciphertext[165]                 =   256'h69c7b273e0f5d06ea4c8880d03064681795bf537c3140b7bf300ffa839d2e5e8;
assign   tb_o_tag_ready[165]                  =   1'b0;
assign   tb_o_tag[165]                        =   tb_o_tag[164];

// CLK no. 166/1240
// *************************************************
assign   tb_i_valid[166]                      =   1'b0;
assign   tb_i_reset[166]                      =   1'b0;
assign   tb_i_sop[166]                        =   1'b0;
assign   tb_i_key_update[166]                 =   1'b0;
assign   tb_i_key[166]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[166]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[166]               =   1'b0;
assign   tb_i_rf_static_encrypt[166]          =   1'b1;
assign   tb_i_clear_fault_flags[166]          =   1'b0;
assign   tb_i_rf_static_aad_length[166]       =   64'h0000000000000100;
assign   tb_i_aad[166]                        =   tb_i_aad[165];
assign   tb_i_rf_static_plaintext_length[166] =   64'h0000000000000280;
assign   tb_i_plaintext[166]                  =   tb_i_plaintext[165];
assign   tb_o_valid[166]                      =   1'b1;
assign   tb_o_sop[166]                        =   1'b0;
assign   tb_o_ciphertext[166]                 =   256'h59c6d418d9f3ac4cbd75e39b25fe803c506469d15f9ba5a9deae5aef075cb038;
assign   tb_o_tag_ready[166]                  =   1'b0;
assign   tb_o_tag[166]                        =   tb_o_tag[165];

// CLK no. 167/1240
// *************************************************
assign   tb_i_valid[167]                      =   1'b0;
assign   tb_i_reset[167]                      =   1'b0;
assign   tb_i_sop[167]                        =   1'b0;
assign   tb_i_key_update[167]                 =   1'b0;
assign   tb_i_key[167]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[167]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[167]               =   1'b0;
assign   tb_i_rf_static_encrypt[167]          =   1'b1;
assign   tb_i_clear_fault_flags[167]          =   1'b0;
assign   tb_i_rf_static_aad_length[167]       =   64'h0000000000000100;
assign   tb_i_aad[167]                        =   tb_i_aad[166];
assign   tb_i_rf_static_plaintext_length[167] =   64'h0000000000000280;
assign   tb_i_plaintext[167]                  =   tb_i_plaintext[166];
assign   tb_o_valid[167]                      =   1'b1;
assign   tb_o_sop[167]                        =   1'b0;
assign   tb_o_ciphertext[167]                 =   256'h80efcf7b82784fb60e2eb6a1b08d8b10;
assign   tb_o_tag_ready[167]                  =   1'b0;
assign   tb_o_tag[167]                        =   tb_o_tag[166];

// CLK no. 168/1240
// *************************************************
assign   tb_i_valid[168]                      =   1'b0;
assign   tb_i_reset[168]                      =   1'b0;
assign   tb_i_sop[168]                        =   1'b0;
assign   tb_i_key_update[168]                 =   1'b0;
assign   tb_i_key[168]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[168]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[168]               =   1'b0;
assign   tb_i_rf_static_encrypt[168]          =   1'b1;
assign   tb_i_clear_fault_flags[168]          =   1'b0;
assign   tb_i_rf_static_aad_length[168]       =   64'h0000000000000100;
assign   tb_i_aad[168]                        =   tb_i_aad[167];
assign   tb_i_rf_static_plaintext_length[168] =   64'h0000000000000280;
assign   tb_i_plaintext[168]                  =   tb_i_plaintext[167];
assign   tb_o_valid[168]                      =   1'b0;
assign   tb_o_sop[168]                        =   1'b0;
assign   tb_o_ciphertext[168]                 =   tb_o_ciphertext[167];
assign   tb_o_tag_ready[168]                  =   1'b0;
assign   tb_o_tag[168]                        =   tb_o_tag[167];

// CLK no. 169/1240
// *************************************************
assign   tb_i_valid[169]                      =   1'b0;
assign   tb_i_reset[169]                      =   1'b0;
assign   tb_i_sop[169]                        =   1'b0;
assign   tb_i_key_update[169]                 =   1'b0;
assign   tb_i_key[169]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[169]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[169]               =   1'b0;
assign   tb_i_rf_static_encrypt[169]          =   1'b1;
assign   tb_i_clear_fault_flags[169]          =   1'b0;
assign   tb_i_rf_static_aad_length[169]       =   64'h0000000000000100;
assign   tb_i_aad[169]                        =   tb_i_aad[168];
assign   tb_i_rf_static_plaintext_length[169] =   64'h0000000000000280;
assign   tb_i_plaintext[169]                  =   tb_i_plaintext[168];
assign   tb_o_valid[169]                      =   1'b0;
assign   tb_o_sop[169]                        =   1'b0;
assign   tb_o_ciphertext[169]                 =   tb_o_ciphertext[168];
assign   tb_o_tag_ready[169]                  =   1'b0;
assign   tb_o_tag[169]                        =   tb_o_tag[168];

// CLK no. 170/1240
// *************************************************
assign   tb_i_valid[170]                      =   1'b0;
assign   tb_i_reset[170]                      =   1'b0;
assign   tb_i_sop[170]                        =   1'b0;
assign   tb_i_key_update[170]                 =   1'b0;
assign   tb_i_key[170]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[170]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[170]               =   1'b0;
assign   tb_i_rf_static_encrypt[170]          =   1'b1;
assign   tb_i_clear_fault_flags[170]          =   1'b0;
assign   tb_i_rf_static_aad_length[170]       =   64'h0000000000000100;
assign   tb_i_aad[170]                        =   tb_i_aad[169];
assign   tb_i_rf_static_plaintext_length[170] =   64'h0000000000000280;
assign   tb_i_plaintext[170]                  =   tb_i_plaintext[169];
assign   tb_o_valid[170]                      =   1'b0;
assign   tb_o_sop[170]                        =   1'b0;
assign   tb_o_ciphertext[170]                 =   tb_o_ciphertext[169];
assign   tb_o_tag_ready[170]                  =   1'b0;
assign   tb_o_tag[170]                        =   tb_o_tag[169];

// CLK no. 171/1240
// *************************************************
assign   tb_i_valid[171]                      =   1'b0;
assign   tb_i_reset[171]                      =   1'b0;
assign   tb_i_sop[171]                        =   1'b0;
assign   tb_i_key_update[171]                 =   1'b0;
assign   tb_i_key[171]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[171]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[171]               =   1'b0;
assign   tb_i_rf_static_encrypt[171]          =   1'b1;
assign   tb_i_clear_fault_flags[171]          =   1'b0;
assign   tb_i_rf_static_aad_length[171]       =   64'h0000000000000100;
assign   tb_i_aad[171]                        =   tb_i_aad[170];
assign   tb_i_rf_static_plaintext_length[171] =   64'h0000000000000280;
assign   tb_i_plaintext[171]                  =   tb_i_plaintext[170];
assign   tb_o_valid[171]                      =   1'b0;
assign   tb_o_sop[171]                        =   1'b0;
assign   tb_o_ciphertext[171]                 =   tb_o_ciphertext[170];
assign   tb_o_tag_ready[171]                  =   1'b0;
assign   tb_o_tag[171]                        =   tb_o_tag[170];

// CLK no. 172/1240
// *************************************************
assign   tb_i_valid[172]                      =   1'b0;
assign   tb_i_reset[172]                      =   1'b0;
assign   tb_i_sop[172]                        =   1'b0;
assign   tb_i_key_update[172]                 =   1'b0;
assign   tb_i_key[172]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[172]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[172]               =   1'b0;
assign   tb_i_rf_static_encrypt[172]          =   1'b1;
assign   tb_i_clear_fault_flags[172]          =   1'b0;
assign   tb_i_rf_static_aad_length[172]       =   64'h0000000000000100;
assign   tb_i_aad[172]                        =   tb_i_aad[171];
assign   tb_i_rf_static_plaintext_length[172] =   64'h0000000000000280;
assign   tb_i_plaintext[172]                  =   tb_i_plaintext[171];
assign   tb_o_valid[172]                      =   1'b0;
assign   tb_o_sop[172]                        =   1'b0;
assign   tb_o_ciphertext[172]                 =   tb_o_ciphertext[171];
assign   tb_o_tag_ready[172]                  =   1'b0;
assign   tb_o_tag[172]                        =   tb_o_tag[171];

// CLK no. 173/1240
// *************************************************
assign   tb_i_valid[173]                      =   1'b0;
assign   tb_i_reset[173]                      =   1'b0;
assign   tb_i_sop[173]                        =   1'b0;
assign   tb_i_key_update[173]                 =   1'b0;
assign   tb_i_key[173]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[173]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[173]               =   1'b0;
assign   tb_i_rf_static_encrypt[173]          =   1'b1;
assign   tb_i_clear_fault_flags[173]          =   1'b0;
assign   tb_i_rf_static_aad_length[173]       =   64'h0000000000000100;
assign   tb_i_aad[173]                        =   tb_i_aad[172];
assign   tb_i_rf_static_plaintext_length[173] =   64'h0000000000000280;
assign   tb_i_plaintext[173]                  =   tb_i_plaintext[172];
assign   tb_o_valid[173]                      =   1'b0;
assign   tb_o_sop[173]                        =   1'b0;
assign   tb_o_ciphertext[173]                 =   tb_o_ciphertext[172];
assign   tb_o_tag_ready[173]                  =   1'b0;
assign   tb_o_tag[173]                        =   tb_o_tag[172];

// CLK no. 174/1240
// *************************************************
assign   tb_i_valid[174]                      =   1'b0;
assign   tb_i_reset[174]                      =   1'b0;
assign   tb_i_sop[174]                        =   1'b0;
assign   tb_i_key_update[174]                 =   1'b0;
assign   tb_i_key[174]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[174]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[174]               =   1'b0;
assign   tb_i_rf_static_encrypt[174]          =   1'b1;
assign   tb_i_clear_fault_flags[174]          =   1'b0;
assign   tb_i_rf_static_aad_length[174]       =   64'h0000000000000100;
assign   tb_i_aad[174]                        =   tb_i_aad[173];
assign   tb_i_rf_static_plaintext_length[174] =   64'h0000000000000280;
assign   tb_i_plaintext[174]                  =   tb_i_plaintext[173];
assign   tb_o_valid[174]                      =   1'b0;
assign   tb_o_sop[174]                        =   1'b0;
assign   tb_o_ciphertext[174]                 =   tb_o_ciphertext[173];
assign   tb_o_tag_ready[174]                  =   1'b0;
assign   tb_o_tag[174]                        =   tb_o_tag[173];

// CLK no. 175/1240
// *************************************************
assign   tb_i_valid[175]                      =   1'b0;
assign   tb_i_reset[175]                      =   1'b0;
assign   tb_i_sop[175]                        =   1'b0;
assign   tb_i_key_update[175]                 =   1'b0;
assign   tb_i_key[175]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[175]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[175]               =   1'b0;
assign   tb_i_rf_static_encrypt[175]          =   1'b1;
assign   tb_i_clear_fault_flags[175]          =   1'b0;
assign   tb_i_rf_static_aad_length[175]       =   64'h0000000000000100;
assign   tb_i_aad[175]                        =   tb_i_aad[174];
assign   tb_i_rf_static_plaintext_length[175] =   64'h0000000000000280;
assign   tb_i_plaintext[175]                  =   tb_i_plaintext[174];
assign   tb_o_valid[175]                      =   1'b0;
assign   tb_o_sop[175]                        =   1'b0;
assign   tb_o_ciphertext[175]                 =   tb_o_ciphertext[174];
assign   tb_o_tag_ready[175]                  =   1'b1;
assign   tb_o_tag[175]                        =   128'h4dd1993f6155018e99352aeeb6194f3d;

// CLK no. 176/1240
// *************************************************
assign   tb_i_valid[176]                      =   1'b0;
assign   tb_i_reset[176]                      =   1'b0;
assign   tb_i_sop[176]                        =   1'b0;
assign   tb_i_key_update[176]                 =   1'b0;
assign   tb_i_key[176]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[176]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[176]               =   1'b0;
assign   tb_i_rf_static_encrypt[176]          =   1'b1;
assign   tb_i_clear_fault_flags[176]          =   1'b0;
assign   tb_i_rf_static_aad_length[176]       =   64'h0000000000000100;
assign   tb_i_aad[176]                        =   tb_i_aad[175];
assign   tb_i_rf_static_plaintext_length[176] =   64'h0000000000000280;
assign   tb_i_plaintext[176]                  =   tb_i_plaintext[175];
assign   tb_o_valid[176]                      =   1'b0;
assign   tb_o_sop[176]                        =   1'b0;
assign   tb_o_ciphertext[176]                 =   tb_o_ciphertext[175];
assign   tb_o_tag_ready[176]                  =   1'b0;
assign   tb_o_tag[176]                        =   tb_o_tag[175];

// CLK no. 177/1240
// *************************************************
assign   tb_i_valid[177]                      =   1'b0;
assign   tb_i_reset[177]                      =   1'b0;
assign   tb_i_sop[177]                        =   1'b0;
assign   tb_i_key_update[177]                 =   1'b0;
assign   tb_i_key[177]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[177]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[177]               =   1'b0;
assign   tb_i_rf_static_encrypt[177]          =   1'b1;
assign   tb_i_clear_fault_flags[177]          =   1'b0;
assign   tb_i_rf_static_aad_length[177]       =   64'h0000000000000100;
assign   tb_i_aad[177]                        =   tb_i_aad[176];
assign   tb_i_rf_static_plaintext_length[177] =   64'h0000000000000280;
assign   tb_i_plaintext[177]                  =   tb_i_plaintext[176];
assign   tb_o_valid[177]                      =   1'b0;
assign   tb_o_sop[177]                        =   1'b0;
assign   tb_o_ciphertext[177]                 =   tb_o_ciphertext[176];
assign   tb_o_tag_ready[177]                  =   1'b0;
assign   tb_o_tag[177]                        =   tb_o_tag[176];

// CLK no. 178/1240
// *************************************************
assign   tb_i_valid[178]                      =   1'b0;
assign   tb_i_reset[178]                      =   1'b0;
assign   tb_i_sop[178]                        =   1'b1;
assign   tb_i_key_update[178]                 =   1'b0;
assign   tb_i_key[178]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[178]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[178]               =   1'b0;
assign   tb_i_rf_static_encrypt[178]          =   1'b1;
assign   tb_i_clear_fault_flags[178]          =   1'b0;
assign   tb_i_rf_static_aad_length[178]       =   64'h0000000000000100;
assign   tb_i_aad[178]                        =   tb_i_aad[177];
assign   tb_i_rf_static_plaintext_length[178] =   64'h0000000000000280;
assign   tb_i_plaintext[178]                  =   tb_i_plaintext[177];
assign   tb_o_valid[178]                      =   1'b0;
assign   tb_o_sop[178]                        =   1'b0;
assign   tb_o_ciphertext[178]                 =   tb_o_ciphertext[177];
assign   tb_o_tag_ready[178]                  =   1'b0;
assign   tb_o_tag[178]                        =   tb_o_tag[177];

// CLK no. 179/1240
// *************************************************
assign   tb_i_valid[179]                      =   1'b1;
assign   tb_i_reset[179]                      =   1'b0;
assign   tb_i_sop[179]                        =   1'b0;
assign   tb_i_key_update[179]                 =   1'b0;
assign   tb_i_key[179]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[179]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[179]               =   1'b0;
assign   tb_i_rf_static_encrypt[179]          =   1'b1;
assign   tb_i_clear_fault_flags[179]          =   1'b0;
assign   tb_i_rf_static_aad_length[179]       =   64'h0000000000000100;
assign   tb_i_aad[179]                        =   256'h1cbffb3b3c7952275f5accf87567dee3c712490db6db5fa317eb373a05b36f9d;
assign   tb_i_rf_static_plaintext_length[179] =   64'h0000000000000280;
assign   tb_i_plaintext[179]                  =   tb_i_plaintext[178];
assign   tb_o_valid[179]                      =   1'b0;
assign   tb_o_sop[179]                        =   1'b0;
assign   tb_o_ciphertext[179]                 =   tb_o_ciphertext[178];
assign   tb_o_tag_ready[179]                  =   1'b0;
assign   tb_o_tag[179]                        =   tb_o_tag[178];

// CLK no. 180/1240
// *************************************************
assign   tb_i_valid[180]                      =   1'b1;
assign   tb_i_reset[180]                      =   1'b0;
assign   tb_i_sop[180]                        =   1'b0;
assign   tb_i_key_update[180]                 =   1'b0;
assign   tb_i_key[180]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[180]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[180]               =   1'b0;
assign   tb_i_rf_static_encrypt[180]          =   1'b1;
assign   tb_i_clear_fault_flags[180]          =   1'b0;
assign   tb_i_rf_static_aad_length[180]       =   64'h0000000000000100;
assign   tb_i_aad[180]                        =   tb_i_aad[179];
assign   tb_i_rf_static_plaintext_length[180] =   64'h0000000000000280;
assign   tb_i_plaintext[180]                  =   256'hfce3021685b85dc839be1afbd9312a587b93dff21223e837c7f6d5636ae05fee;
assign   tb_o_valid[180]                      =   1'b0;
assign   tb_o_sop[180]                        =   1'b0;
assign   tb_o_ciphertext[180]                 =   tb_o_ciphertext[179];
assign   tb_o_tag_ready[180]                  =   1'b0;
assign   tb_o_tag[180]                        =   tb_o_tag[179];

// CLK no. 181/1240
// *************************************************
assign   tb_i_valid[181]                      =   1'b1;
assign   tb_i_reset[181]                      =   1'b0;
assign   tb_i_sop[181]                        =   1'b0;
assign   tb_i_key_update[181]                 =   1'b0;
assign   tb_i_key[181]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[181]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[181]               =   1'b0;
assign   tb_i_rf_static_encrypt[181]          =   1'b1;
assign   tb_i_clear_fault_flags[181]          =   1'b0;
assign   tb_i_rf_static_aad_length[181]       =   64'h0000000000000100;
assign   tb_i_aad[181]                        =   tb_i_aad[180];
assign   tb_i_rf_static_plaintext_length[181] =   64'h0000000000000280;
assign   tb_i_plaintext[181]                  =   256'h6ea82714ed7f30046729f3def1850bb32ad667d9324e21103d5f069944128f13;
assign   tb_o_valid[181]                      =   1'b0;
assign   tb_o_sop[181]                        =   1'b0;
assign   tb_o_ciphertext[181]                 =   tb_o_ciphertext[180];
assign   tb_o_tag_ready[181]                  =   1'b0;
assign   tb_o_tag[181]                        =   tb_o_tag[180];

// CLK no. 182/1240
// *************************************************
assign   tb_i_valid[182]                      =   1'b1;
assign   tb_i_reset[182]                      =   1'b0;
assign   tb_i_sop[182]                        =   1'b0;
assign   tb_i_key_update[182]                 =   1'b0;
assign   tb_i_key[182]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[182]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[182]               =   1'b0;
assign   tb_i_rf_static_encrypt[182]          =   1'b1;
assign   tb_i_clear_fault_flags[182]          =   1'b0;
assign   tb_i_rf_static_aad_length[182]       =   64'h0000000000000100;
assign   tb_i_aad[182]                        =   tb_i_aad[181];
assign   tb_i_rf_static_plaintext_length[182] =   64'h0000000000000280;
assign   tb_i_plaintext[182]                  =   256'h12bca566310979cdcec19f88dcefa24b;
assign   tb_o_valid[182]                      =   1'b0;
assign   tb_o_sop[182]                        =   1'b0;
assign   tb_o_ciphertext[182]                 =   tb_o_ciphertext[181];
assign   tb_o_tag_ready[182]                  =   1'b0;
assign   tb_o_tag[182]                        =   tb_o_tag[181];

// CLK no. 183/1240
// *************************************************
assign   tb_i_valid[183]                      =   1'b0;
assign   tb_i_reset[183]                      =   1'b0;
assign   tb_i_sop[183]                        =   1'b0;
assign   tb_i_key_update[183]                 =   1'b0;
assign   tb_i_key[183]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[183]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[183]               =   1'b0;
assign   tb_i_rf_static_encrypt[183]          =   1'b1;
assign   tb_i_clear_fault_flags[183]          =   1'b0;
assign   tb_i_rf_static_aad_length[183]       =   64'h0000000000000100;
assign   tb_i_aad[183]                        =   tb_i_aad[182];
assign   tb_i_rf_static_plaintext_length[183] =   64'h0000000000000280;
assign   tb_i_plaintext[183]                  =   tb_i_plaintext[182];
assign   tb_o_valid[183]                      =   1'b0;
assign   tb_o_sop[183]                        =   1'b0;
assign   tb_o_ciphertext[183]                 =   tb_o_ciphertext[182];
assign   tb_o_tag_ready[183]                  =   1'b0;
assign   tb_o_tag[183]                        =   tb_o_tag[182];

// CLK no. 184/1240
// *************************************************
assign   tb_i_valid[184]                      =   1'b0;
assign   tb_i_reset[184]                      =   1'b0;
assign   tb_i_sop[184]                        =   1'b0;
assign   tb_i_key_update[184]                 =   1'b0;
assign   tb_i_key[184]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[184]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[184]               =   1'b0;
assign   tb_i_rf_static_encrypt[184]          =   1'b1;
assign   tb_i_clear_fault_flags[184]          =   1'b0;
assign   tb_i_rf_static_aad_length[184]       =   64'h0000000000000100;
assign   tb_i_aad[184]                        =   tb_i_aad[183];
assign   tb_i_rf_static_plaintext_length[184] =   64'h0000000000000280;
assign   tb_i_plaintext[184]                  =   tb_i_plaintext[183];
assign   tb_o_valid[184]                      =   1'b0;
assign   tb_o_sop[184]                        =   1'b0;
assign   tb_o_ciphertext[184]                 =   tb_o_ciphertext[183];
assign   tb_o_tag_ready[184]                  =   1'b0;
assign   tb_o_tag[184]                        =   tb_o_tag[183];

// CLK no. 185/1240
// *************************************************
assign   tb_i_valid[185]                      =   1'b0;
assign   tb_i_reset[185]                      =   1'b0;
assign   tb_i_sop[185]                        =   1'b0;
assign   tb_i_key_update[185]                 =   1'b0;
assign   tb_i_key[185]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[185]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[185]               =   1'b0;
assign   tb_i_rf_static_encrypt[185]          =   1'b1;
assign   tb_i_clear_fault_flags[185]          =   1'b0;
assign   tb_i_rf_static_aad_length[185]       =   64'h0000000000000100;
assign   tb_i_aad[185]                        =   tb_i_aad[184];
assign   tb_i_rf_static_plaintext_length[185] =   64'h0000000000000280;
assign   tb_i_plaintext[185]                  =   tb_i_plaintext[184];
assign   tb_o_valid[185]                      =   1'b0;
assign   tb_o_sop[185]                        =   1'b0;
assign   tb_o_ciphertext[185]                 =   tb_o_ciphertext[184];
assign   tb_o_tag_ready[185]                  =   1'b0;
assign   tb_o_tag[185]                        =   tb_o_tag[184];

// CLK no. 186/1240
// *************************************************
assign   tb_i_valid[186]                      =   1'b0;
assign   tb_i_reset[186]                      =   1'b0;
assign   tb_i_sop[186]                        =   1'b0;
assign   tb_i_key_update[186]                 =   1'b0;
assign   tb_i_key[186]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[186]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[186]               =   1'b0;
assign   tb_i_rf_static_encrypt[186]          =   1'b1;
assign   tb_i_clear_fault_flags[186]          =   1'b0;
assign   tb_i_rf_static_aad_length[186]       =   64'h0000000000000100;
assign   tb_i_aad[186]                        =   tb_i_aad[185];
assign   tb_i_rf_static_plaintext_length[186] =   64'h0000000000000280;
assign   tb_i_plaintext[186]                  =   tb_i_plaintext[185];
assign   tb_o_valid[186]                      =   1'b0;
assign   tb_o_sop[186]                        =   1'b0;
assign   tb_o_ciphertext[186]                 =   tb_o_ciphertext[185];
assign   tb_o_tag_ready[186]                  =   1'b0;
assign   tb_o_tag[186]                        =   tb_o_tag[185];

// CLK no. 187/1240
// *************************************************
assign   tb_i_valid[187]                      =   1'b0;
assign   tb_i_reset[187]                      =   1'b0;
assign   tb_i_sop[187]                        =   1'b0;
assign   tb_i_key_update[187]                 =   1'b0;
assign   tb_i_key[187]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[187]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[187]               =   1'b0;
assign   tb_i_rf_static_encrypt[187]          =   1'b1;
assign   tb_i_clear_fault_flags[187]          =   1'b0;
assign   tb_i_rf_static_aad_length[187]       =   64'h0000000000000100;
assign   tb_i_aad[187]                        =   tb_i_aad[186];
assign   tb_i_rf_static_plaintext_length[187] =   64'h0000000000000280;
assign   tb_i_plaintext[187]                  =   tb_i_plaintext[186];
assign   tb_o_valid[187]                      =   1'b0;
assign   tb_o_sop[187]                        =   1'b0;
assign   tb_o_ciphertext[187]                 =   tb_o_ciphertext[186];
assign   tb_o_tag_ready[187]                  =   1'b0;
assign   tb_o_tag[187]                        =   tb_o_tag[186];

// CLK no. 188/1240
// *************************************************
assign   tb_i_valid[188]                      =   1'b0;
assign   tb_i_reset[188]                      =   1'b0;
assign   tb_i_sop[188]                        =   1'b0;
assign   tb_i_key_update[188]                 =   1'b0;
assign   tb_i_key[188]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[188]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[188]               =   1'b0;
assign   tb_i_rf_static_encrypt[188]          =   1'b1;
assign   tb_i_clear_fault_flags[188]          =   1'b0;
assign   tb_i_rf_static_aad_length[188]       =   64'h0000000000000100;
assign   tb_i_aad[188]                        =   tb_i_aad[187];
assign   tb_i_rf_static_plaintext_length[188] =   64'h0000000000000280;
assign   tb_i_plaintext[188]                  =   tb_i_plaintext[187];
assign   tb_o_valid[188]                      =   1'b0;
assign   tb_o_sop[188]                        =   1'b0;
assign   tb_o_ciphertext[188]                 =   tb_o_ciphertext[187];
assign   tb_o_tag_ready[188]                  =   1'b0;
assign   tb_o_tag[188]                        =   tb_o_tag[187];

// CLK no. 189/1240
// *************************************************
assign   tb_i_valid[189]                      =   1'b0;
assign   tb_i_reset[189]                      =   1'b0;
assign   tb_i_sop[189]                        =   1'b0;
assign   tb_i_key_update[189]                 =   1'b0;
assign   tb_i_key[189]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[189]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[189]               =   1'b0;
assign   tb_i_rf_static_encrypt[189]          =   1'b1;
assign   tb_i_clear_fault_flags[189]          =   1'b0;
assign   tb_i_rf_static_aad_length[189]       =   64'h0000000000000100;
assign   tb_i_aad[189]                        =   tb_i_aad[188];
assign   tb_i_rf_static_plaintext_length[189] =   64'h0000000000000280;
assign   tb_i_plaintext[189]                  =   tb_i_plaintext[188];
assign   tb_o_valid[189]                      =   1'b0;
assign   tb_o_sop[189]                        =   1'b0;
assign   tb_o_ciphertext[189]                 =   tb_o_ciphertext[188];
assign   tb_o_tag_ready[189]                  =   1'b0;
assign   tb_o_tag[189]                        =   tb_o_tag[188];

// CLK no. 190/1240
// *************************************************
assign   tb_i_valid[190]                      =   1'b0;
assign   tb_i_reset[190]                      =   1'b0;
assign   tb_i_sop[190]                        =   1'b0;
assign   tb_i_key_update[190]                 =   1'b0;
assign   tb_i_key[190]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[190]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[190]               =   1'b0;
assign   tb_i_rf_static_encrypt[190]          =   1'b1;
assign   tb_i_clear_fault_flags[190]          =   1'b0;
assign   tb_i_rf_static_aad_length[190]       =   64'h0000000000000100;
assign   tb_i_aad[190]                        =   tb_i_aad[189];
assign   tb_i_rf_static_plaintext_length[190] =   64'h0000000000000280;
assign   tb_i_plaintext[190]                  =   tb_i_plaintext[189];
assign   tb_o_valid[190]                      =   1'b0;
assign   tb_o_sop[190]                        =   1'b0;
assign   tb_o_ciphertext[190]                 =   tb_o_ciphertext[189];
assign   tb_o_tag_ready[190]                  =   1'b0;
assign   tb_o_tag[190]                        =   tb_o_tag[189];

// CLK no. 191/1240
// *************************************************
assign   tb_i_valid[191]                      =   1'b0;
assign   tb_i_reset[191]                      =   1'b0;
assign   tb_i_sop[191]                        =   1'b0;
assign   tb_i_key_update[191]                 =   1'b0;
assign   tb_i_key[191]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[191]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[191]               =   1'b0;
assign   tb_i_rf_static_encrypt[191]          =   1'b1;
assign   tb_i_clear_fault_flags[191]          =   1'b0;
assign   tb_i_rf_static_aad_length[191]       =   64'h0000000000000100;
assign   tb_i_aad[191]                        =   tb_i_aad[190];
assign   tb_i_rf_static_plaintext_length[191] =   64'h0000000000000280;
assign   tb_i_plaintext[191]                  =   tb_i_plaintext[190];
assign   tb_o_valid[191]                      =   1'b0;
assign   tb_o_sop[191]                        =   1'b0;
assign   tb_o_ciphertext[191]                 =   tb_o_ciphertext[190];
assign   tb_o_tag_ready[191]                  =   1'b0;
assign   tb_o_tag[191]                        =   tb_o_tag[190];

// CLK no. 192/1240
// *************************************************
assign   tb_i_valid[192]                      =   1'b0;
assign   tb_i_reset[192]                      =   1'b0;
assign   tb_i_sop[192]                        =   1'b0;
assign   tb_i_key_update[192]                 =   1'b0;
assign   tb_i_key[192]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[192]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[192]               =   1'b0;
assign   tb_i_rf_static_encrypt[192]          =   1'b1;
assign   tb_i_clear_fault_flags[192]          =   1'b0;
assign   tb_i_rf_static_aad_length[192]       =   64'h0000000000000100;
assign   tb_i_aad[192]                        =   tb_i_aad[191];
assign   tb_i_rf_static_plaintext_length[192] =   64'h0000000000000280;
assign   tb_i_plaintext[192]                  =   tb_i_plaintext[191];
assign   tb_o_valid[192]                      =   1'b0;
assign   tb_o_sop[192]                        =   1'b0;
assign   tb_o_ciphertext[192]                 =   tb_o_ciphertext[191];
assign   tb_o_tag_ready[192]                  =   1'b0;
assign   tb_o_tag[192]                        =   tb_o_tag[191];

// CLK no. 193/1240
// *************************************************
assign   tb_i_valid[193]                      =   1'b0;
assign   tb_i_reset[193]                      =   1'b0;
assign   tb_i_sop[193]                        =   1'b0;
assign   tb_i_key_update[193]                 =   1'b0;
assign   tb_i_key[193]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[193]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[193]               =   1'b0;
assign   tb_i_rf_static_encrypt[193]          =   1'b1;
assign   tb_i_clear_fault_flags[193]          =   1'b0;
assign   tb_i_rf_static_aad_length[193]       =   64'h0000000000000100;
assign   tb_i_aad[193]                        =   tb_i_aad[192];
assign   tb_i_rf_static_plaintext_length[193] =   64'h0000000000000280;
assign   tb_i_plaintext[193]                  =   tb_i_plaintext[192];
assign   tb_o_valid[193]                      =   1'b0;
assign   tb_o_sop[193]                        =   1'b0;
assign   tb_o_ciphertext[193]                 =   tb_o_ciphertext[192];
assign   tb_o_tag_ready[193]                  =   1'b0;
assign   tb_o_tag[193]                        =   tb_o_tag[192];

// CLK no. 194/1240
// *************************************************
assign   tb_i_valid[194]                      =   1'b0;
assign   tb_i_reset[194]                      =   1'b0;
assign   tb_i_sop[194]                        =   1'b0;
assign   tb_i_key_update[194]                 =   1'b0;
assign   tb_i_key[194]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[194]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[194]               =   1'b0;
assign   tb_i_rf_static_encrypt[194]          =   1'b1;
assign   tb_i_clear_fault_flags[194]          =   1'b0;
assign   tb_i_rf_static_aad_length[194]       =   64'h0000000000000100;
assign   tb_i_aad[194]                        =   tb_i_aad[193];
assign   tb_i_rf_static_plaintext_length[194] =   64'h0000000000000280;
assign   tb_i_plaintext[194]                  =   tb_i_plaintext[193];
assign   tb_o_valid[194]                      =   1'b0;
assign   tb_o_sop[194]                        =   1'b0;
assign   tb_o_ciphertext[194]                 =   tb_o_ciphertext[193];
assign   tb_o_tag_ready[194]                  =   1'b0;
assign   tb_o_tag[194]                        =   tb_o_tag[193];

// CLK no. 195/1240
// *************************************************
assign   tb_i_valid[195]                      =   1'b0;
assign   tb_i_reset[195]                      =   1'b0;
assign   tb_i_sop[195]                        =   1'b0;
assign   tb_i_key_update[195]                 =   1'b0;
assign   tb_i_key[195]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[195]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[195]               =   1'b0;
assign   tb_i_rf_static_encrypt[195]          =   1'b1;
assign   tb_i_clear_fault_flags[195]          =   1'b0;
assign   tb_i_rf_static_aad_length[195]       =   64'h0000000000000100;
assign   tb_i_aad[195]                        =   tb_i_aad[194];
assign   tb_i_rf_static_plaintext_length[195] =   64'h0000000000000280;
assign   tb_i_plaintext[195]                  =   tb_i_plaintext[194];
assign   tb_o_valid[195]                      =   1'b0;
assign   tb_o_sop[195]                        =   1'b0;
assign   tb_o_ciphertext[195]                 =   tb_o_ciphertext[194];
assign   tb_o_tag_ready[195]                  =   1'b0;
assign   tb_o_tag[195]                        =   tb_o_tag[194];

// CLK no. 196/1240
// *************************************************
assign   tb_i_valid[196]                      =   1'b0;
assign   tb_i_reset[196]                      =   1'b0;
assign   tb_i_sop[196]                        =   1'b0;
assign   tb_i_key_update[196]                 =   1'b0;
assign   tb_i_key[196]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[196]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[196]               =   1'b0;
assign   tb_i_rf_static_encrypt[196]          =   1'b1;
assign   tb_i_clear_fault_flags[196]          =   1'b0;
assign   tb_i_rf_static_aad_length[196]       =   64'h0000000000000100;
assign   tb_i_aad[196]                        =   tb_i_aad[195];
assign   tb_i_rf_static_plaintext_length[196] =   64'h0000000000000280;
assign   tb_i_plaintext[196]                  =   tb_i_plaintext[195];
assign   tb_o_valid[196]                      =   1'b0;
assign   tb_o_sop[196]                        =   1'b0;
assign   tb_o_ciphertext[196]                 =   tb_o_ciphertext[195];
assign   tb_o_tag_ready[196]                  =   1'b0;
assign   tb_o_tag[196]                        =   tb_o_tag[195];

// CLK no. 197/1240
// *************************************************
assign   tb_i_valid[197]                      =   1'b0;
assign   tb_i_reset[197]                      =   1'b0;
assign   tb_i_sop[197]                        =   1'b0;
assign   tb_i_key_update[197]                 =   1'b0;
assign   tb_i_key[197]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[197]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[197]               =   1'b0;
assign   tb_i_rf_static_encrypt[197]          =   1'b1;
assign   tb_i_clear_fault_flags[197]          =   1'b0;
assign   tb_i_rf_static_aad_length[197]       =   64'h0000000000000100;
assign   tb_i_aad[197]                        =   tb_i_aad[196];
assign   tb_i_rf_static_plaintext_length[197] =   64'h0000000000000280;
assign   tb_i_plaintext[197]                  =   tb_i_plaintext[196];
assign   tb_o_valid[197]                      =   1'b0;
assign   tb_o_sop[197]                        =   1'b0;
assign   tb_o_ciphertext[197]                 =   tb_o_ciphertext[196];
assign   tb_o_tag_ready[197]                  =   1'b0;
assign   tb_o_tag[197]                        =   tb_o_tag[196];

// CLK no. 198/1240
// *************************************************
assign   tb_i_valid[198]                      =   1'b0;
assign   tb_i_reset[198]                      =   1'b0;
assign   tb_i_sop[198]                        =   1'b0;
assign   tb_i_key_update[198]                 =   1'b0;
assign   tb_i_key[198]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[198]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[198]               =   1'b0;
assign   tb_i_rf_static_encrypt[198]          =   1'b1;
assign   tb_i_clear_fault_flags[198]          =   1'b0;
assign   tb_i_rf_static_aad_length[198]       =   64'h0000000000000100;
assign   tb_i_aad[198]                        =   tb_i_aad[197];
assign   tb_i_rf_static_plaintext_length[198] =   64'h0000000000000280;
assign   tb_i_plaintext[198]                  =   tb_i_plaintext[197];
assign   tb_o_valid[198]                      =   1'b0;
assign   tb_o_sop[198]                        =   1'b0;
assign   tb_o_ciphertext[198]                 =   tb_o_ciphertext[197];
assign   tb_o_tag_ready[198]                  =   1'b0;
assign   tb_o_tag[198]                        =   tb_o_tag[197];

// CLK no. 199/1240
// *************************************************
assign   tb_i_valid[199]                      =   1'b0;
assign   tb_i_reset[199]                      =   1'b0;
assign   tb_i_sop[199]                        =   1'b0;
assign   tb_i_key_update[199]                 =   1'b0;
assign   tb_i_key[199]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[199]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[199]               =   1'b0;
assign   tb_i_rf_static_encrypt[199]          =   1'b1;
assign   tb_i_clear_fault_flags[199]          =   1'b0;
assign   tb_i_rf_static_aad_length[199]       =   64'h0000000000000100;
assign   tb_i_aad[199]                        =   tb_i_aad[198];
assign   tb_i_rf_static_plaintext_length[199] =   64'h0000000000000280;
assign   tb_i_plaintext[199]                  =   tb_i_plaintext[198];
assign   tb_o_valid[199]                      =   1'b0;
assign   tb_o_sop[199]                        =   1'b0;
assign   tb_o_ciphertext[199]                 =   tb_o_ciphertext[198];
assign   tb_o_tag_ready[199]                  =   1'b0;
assign   tb_o_tag[199]                        =   tb_o_tag[198];

// CLK no. 200/1240
// *************************************************
assign   tb_i_valid[200]                      =   1'b0;
assign   tb_i_reset[200]                      =   1'b0;
assign   tb_i_sop[200]                        =   1'b0;
assign   tb_i_key_update[200]                 =   1'b0;
assign   tb_i_key[200]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[200]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[200]               =   1'b0;
assign   tb_i_rf_static_encrypt[200]          =   1'b1;
assign   tb_i_clear_fault_flags[200]          =   1'b0;
assign   tb_i_rf_static_aad_length[200]       =   64'h0000000000000100;
assign   tb_i_aad[200]                        =   tb_i_aad[199];
assign   tb_i_rf_static_plaintext_length[200] =   64'h0000000000000280;
assign   tb_i_plaintext[200]                  =   tb_i_plaintext[199];
assign   tb_o_valid[200]                      =   1'b0;
assign   tb_o_sop[200]                        =   1'b0;
assign   tb_o_ciphertext[200]                 =   tb_o_ciphertext[199];
assign   tb_o_tag_ready[200]                  =   1'b0;
assign   tb_o_tag[200]                        =   tb_o_tag[199];

// CLK no. 201/1240
// *************************************************
assign   tb_i_valid[201]                      =   1'b0;
assign   tb_i_reset[201]                      =   1'b0;
assign   tb_i_sop[201]                        =   1'b0;
assign   tb_i_key_update[201]                 =   1'b0;
assign   tb_i_key[201]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[201]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[201]               =   1'b0;
assign   tb_i_rf_static_encrypt[201]          =   1'b1;
assign   tb_i_clear_fault_flags[201]          =   1'b0;
assign   tb_i_rf_static_aad_length[201]       =   64'h0000000000000100;
assign   tb_i_aad[201]                        =   tb_i_aad[200];
assign   tb_i_rf_static_plaintext_length[201] =   64'h0000000000000280;
assign   tb_i_plaintext[201]                  =   tb_i_plaintext[200];
assign   tb_o_valid[201]                      =   1'b0;
assign   tb_o_sop[201]                        =   1'b0;
assign   tb_o_ciphertext[201]                 =   tb_o_ciphertext[200];
assign   tb_o_tag_ready[201]                  =   1'b0;
assign   tb_o_tag[201]                        =   tb_o_tag[200];

// CLK no. 202/1240
// *************************************************
assign   tb_i_valid[202]                      =   1'b0;
assign   tb_i_reset[202]                      =   1'b0;
assign   tb_i_sop[202]                        =   1'b0;
assign   tb_i_key_update[202]                 =   1'b0;
assign   tb_i_key[202]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[202]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[202]               =   1'b0;
assign   tb_i_rf_static_encrypt[202]          =   1'b1;
assign   tb_i_clear_fault_flags[202]          =   1'b0;
assign   tb_i_rf_static_aad_length[202]       =   64'h0000000000000100;
assign   tb_i_aad[202]                        =   tb_i_aad[201];
assign   tb_i_rf_static_plaintext_length[202] =   64'h0000000000000280;
assign   tb_i_plaintext[202]                  =   tb_i_plaintext[201];
assign   tb_o_valid[202]                      =   1'b0;
assign   tb_o_sop[202]                        =   1'b0;
assign   tb_o_ciphertext[202]                 =   tb_o_ciphertext[201];
assign   tb_o_tag_ready[202]                  =   1'b0;
assign   tb_o_tag[202]                        =   tb_o_tag[201];

// CLK no. 203/1240
// *************************************************
assign   tb_i_valid[203]                      =   1'b0;
assign   tb_i_reset[203]                      =   1'b0;
assign   tb_i_sop[203]                        =   1'b0;
assign   tb_i_key_update[203]                 =   1'b0;
assign   tb_i_key[203]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[203]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[203]               =   1'b0;
assign   tb_i_rf_static_encrypt[203]          =   1'b1;
assign   tb_i_clear_fault_flags[203]          =   1'b0;
assign   tb_i_rf_static_aad_length[203]       =   64'h0000000000000100;
assign   tb_i_aad[203]                        =   tb_i_aad[202];
assign   tb_i_rf_static_plaintext_length[203] =   64'h0000000000000280;
assign   tb_i_plaintext[203]                  =   tb_i_plaintext[202];
assign   tb_o_valid[203]                      =   1'b0;
assign   tb_o_sop[203]                        =   1'b0;
assign   tb_o_ciphertext[203]                 =   tb_o_ciphertext[202];
assign   tb_o_tag_ready[203]                  =   1'b0;
assign   tb_o_tag[203]                        =   tb_o_tag[202];

// CLK no. 204/1240
// *************************************************
assign   tb_i_valid[204]                      =   1'b0;
assign   tb_i_reset[204]                      =   1'b0;
assign   tb_i_sop[204]                        =   1'b0;
assign   tb_i_key_update[204]                 =   1'b0;
assign   tb_i_key[204]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[204]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[204]               =   1'b0;
assign   tb_i_rf_static_encrypt[204]          =   1'b1;
assign   tb_i_clear_fault_flags[204]          =   1'b0;
assign   tb_i_rf_static_aad_length[204]       =   64'h0000000000000100;
assign   tb_i_aad[204]                        =   tb_i_aad[203];
assign   tb_i_rf_static_plaintext_length[204] =   64'h0000000000000280;
assign   tb_i_plaintext[204]                  =   tb_i_plaintext[203];
assign   tb_o_valid[204]                      =   1'b0;
assign   tb_o_sop[204]                        =   1'b0;
assign   tb_o_ciphertext[204]                 =   tb_o_ciphertext[203];
assign   tb_o_tag_ready[204]                  =   1'b0;
assign   tb_o_tag[204]                        =   tb_o_tag[203];

// CLK no. 205/1240
// *************************************************
assign   tb_i_valid[205]                      =   1'b0;
assign   tb_i_reset[205]                      =   1'b0;
assign   tb_i_sop[205]                        =   1'b0;
assign   tb_i_key_update[205]                 =   1'b0;
assign   tb_i_key[205]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[205]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[205]               =   1'b0;
assign   tb_i_rf_static_encrypt[205]          =   1'b1;
assign   tb_i_clear_fault_flags[205]          =   1'b0;
assign   tb_i_rf_static_aad_length[205]       =   64'h0000000000000100;
assign   tb_i_aad[205]                        =   tb_i_aad[204];
assign   tb_i_rf_static_plaintext_length[205] =   64'h0000000000000280;
assign   tb_i_plaintext[205]                  =   tb_i_plaintext[204];
assign   tb_o_valid[205]                      =   1'b0;
assign   tb_o_sop[205]                        =   1'b0;
assign   tb_o_ciphertext[205]                 =   tb_o_ciphertext[204];
assign   tb_o_tag_ready[205]                  =   1'b0;
assign   tb_o_tag[205]                        =   tb_o_tag[204];

// CLK no. 206/1240
// *************************************************
assign   tb_i_valid[206]                      =   1'b0;
assign   tb_i_reset[206]                      =   1'b0;
assign   tb_i_sop[206]                        =   1'b0;
assign   tb_i_key_update[206]                 =   1'b0;
assign   tb_i_key[206]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[206]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[206]               =   1'b0;
assign   tb_i_rf_static_encrypt[206]          =   1'b1;
assign   tb_i_clear_fault_flags[206]          =   1'b0;
assign   tb_i_rf_static_aad_length[206]       =   64'h0000000000000100;
assign   tb_i_aad[206]                        =   tb_i_aad[205];
assign   tb_i_rf_static_plaintext_length[206] =   64'h0000000000000280;
assign   tb_i_plaintext[206]                  =   tb_i_plaintext[205];
assign   tb_o_valid[206]                      =   1'b0;
assign   tb_o_sop[206]                        =   1'b0;
assign   tb_o_ciphertext[206]                 =   tb_o_ciphertext[205];
assign   tb_o_tag_ready[206]                  =   1'b0;
assign   tb_o_tag[206]                        =   tb_o_tag[205];

// CLK no. 207/1240
// *************************************************
assign   tb_i_valid[207]                      =   1'b0;
assign   tb_i_reset[207]                      =   1'b0;
assign   tb_i_sop[207]                        =   1'b0;
assign   tb_i_key_update[207]                 =   1'b0;
assign   tb_i_key[207]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[207]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[207]               =   1'b0;
assign   tb_i_rf_static_encrypt[207]          =   1'b1;
assign   tb_i_clear_fault_flags[207]          =   1'b0;
assign   tb_i_rf_static_aad_length[207]       =   64'h0000000000000100;
assign   tb_i_aad[207]                        =   tb_i_aad[206];
assign   tb_i_rf_static_plaintext_length[207] =   64'h0000000000000280;
assign   tb_i_plaintext[207]                  =   tb_i_plaintext[206];
assign   tb_o_valid[207]                      =   1'b0;
assign   tb_o_sop[207]                        =   1'b0;
assign   tb_o_ciphertext[207]                 =   tb_o_ciphertext[206];
assign   tb_o_tag_ready[207]                  =   1'b0;
assign   tb_o_tag[207]                        =   tb_o_tag[206];

// CLK no. 208/1240
// *************************************************
assign   tb_i_valid[208]                      =   1'b0;
assign   tb_i_reset[208]                      =   1'b0;
assign   tb_i_sop[208]                        =   1'b0;
assign   tb_i_key_update[208]                 =   1'b0;
assign   tb_i_key[208]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[208]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[208]               =   1'b0;
assign   tb_i_rf_static_encrypt[208]          =   1'b1;
assign   tb_i_clear_fault_flags[208]          =   1'b0;
assign   tb_i_rf_static_aad_length[208]       =   64'h0000000000000100;
assign   tb_i_aad[208]                        =   tb_i_aad[207];
assign   tb_i_rf_static_plaintext_length[208] =   64'h0000000000000280;
assign   tb_i_plaintext[208]                  =   tb_i_plaintext[207];
assign   tb_o_valid[208]                      =   1'b0;
assign   tb_o_sop[208]                        =   1'b0;
assign   tb_o_ciphertext[208]                 =   tb_o_ciphertext[207];
assign   tb_o_tag_ready[208]                  =   1'b0;
assign   tb_o_tag[208]                        =   tb_o_tag[207];

// CLK no. 209/1240
// *************************************************
assign   tb_i_valid[209]                      =   1'b0;
assign   tb_i_reset[209]                      =   1'b0;
assign   tb_i_sop[209]                        =   1'b0;
assign   tb_i_key_update[209]                 =   1'b0;
assign   tb_i_key[209]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[209]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[209]               =   1'b0;
assign   tb_i_rf_static_encrypt[209]          =   1'b1;
assign   tb_i_clear_fault_flags[209]          =   1'b0;
assign   tb_i_rf_static_aad_length[209]       =   64'h0000000000000100;
assign   tb_i_aad[209]                        =   tb_i_aad[208];
assign   tb_i_rf_static_plaintext_length[209] =   64'h0000000000000280;
assign   tb_i_plaintext[209]                  =   tb_i_plaintext[208];
assign   tb_o_valid[209]                      =   1'b0;
assign   tb_o_sop[209]                        =   1'b0;
assign   tb_o_ciphertext[209]                 =   tb_o_ciphertext[208];
assign   tb_o_tag_ready[209]                  =   1'b0;
assign   tb_o_tag[209]                        =   tb_o_tag[208];

// CLK no. 210/1240
// *************************************************
assign   tb_i_valid[210]                      =   1'b0;
assign   tb_i_reset[210]                      =   1'b0;
assign   tb_i_sop[210]                        =   1'b0;
assign   tb_i_key_update[210]                 =   1'b0;
assign   tb_i_key[210]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[210]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[210]               =   1'b0;
assign   tb_i_rf_static_encrypt[210]          =   1'b1;
assign   tb_i_clear_fault_flags[210]          =   1'b0;
assign   tb_i_rf_static_aad_length[210]       =   64'h0000000000000100;
assign   tb_i_aad[210]                        =   tb_i_aad[209];
assign   tb_i_rf_static_plaintext_length[210] =   64'h0000000000000280;
assign   tb_i_plaintext[210]                  =   tb_i_plaintext[209];
assign   tb_o_valid[210]                      =   1'b0;
assign   tb_o_sop[210]                        =   1'b0;
assign   tb_o_ciphertext[210]                 =   tb_o_ciphertext[209];
assign   tb_o_tag_ready[210]                  =   1'b0;
assign   tb_o_tag[210]                        =   tb_o_tag[209];

// CLK no. 211/1240
// *************************************************
assign   tb_i_valid[211]                      =   1'b0;
assign   tb_i_reset[211]                      =   1'b0;
assign   tb_i_sop[211]                        =   1'b0;
assign   tb_i_key_update[211]                 =   1'b0;
assign   tb_i_key[211]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[211]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[211]               =   1'b0;
assign   tb_i_rf_static_encrypt[211]          =   1'b1;
assign   tb_i_clear_fault_flags[211]          =   1'b0;
assign   tb_i_rf_static_aad_length[211]       =   64'h0000000000000100;
assign   tb_i_aad[211]                        =   tb_i_aad[210];
assign   tb_i_rf_static_plaintext_length[211] =   64'h0000000000000280;
assign   tb_i_plaintext[211]                  =   tb_i_plaintext[210];
assign   tb_o_valid[211]                      =   1'b0;
assign   tb_o_sop[211]                        =   1'b0;
assign   tb_o_ciphertext[211]                 =   tb_o_ciphertext[210];
assign   tb_o_tag_ready[211]                  =   1'b0;
assign   tb_o_tag[211]                        =   tb_o_tag[210];

// CLK no. 212/1240
// *************************************************
assign   tb_i_valid[212]                      =   1'b0;
assign   tb_i_reset[212]                      =   1'b0;
assign   tb_i_sop[212]                        =   1'b0;
assign   tb_i_key_update[212]                 =   1'b0;
assign   tb_i_key[212]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[212]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[212]               =   1'b0;
assign   tb_i_rf_static_encrypt[212]          =   1'b1;
assign   tb_i_clear_fault_flags[212]          =   1'b0;
assign   tb_i_rf_static_aad_length[212]       =   64'h0000000000000100;
assign   tb_i_aad[212]                        =   tb_i_aad[211];
assign   tb_i_rf_static_plaintext_length[212] =   64'h0000000000000280;
assign   tb_i_plaintext[212]                  =   tb_i_plaintext[211];
assign   tb_o_valid[212]                      =   1'b0;
assign   tb_o_sop[212]                        =   1'b0;
assign   tb_o_ciphertext[212]                 =   tb_o_ciphertext[211];
assign   tb_o_tag_ready[212]                  =   1'b0;
assign   tb_o_tag[212]                        =   tb_o_tag[211];

// CLK no. 213/1240
// *************************************************
assign   tb_i_valid[213]                      =   1'b0;
assign   tb_i_reset[213]                      =   1'b0;
assign   tb_i_sop[213]                        =   1'b0;
assign   tb_i_key_update[213]                 =   1'b0;
assign   tb_i_key[213]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[213]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[213]               =   1'b0;
assign   tb_i_rf_static_encrypt[213]          =   1'b1;
assign   tb_i_clear_fault_flags[213]          =   1'b0;
assign   tb_i_rf_static_aad_length[213]       =   64'h0000000000000100;
assign   tb_i_aad[213]                        =   tb_i_aad[212];
assign   tb_i_rf_static_plaintext_length[213] =   64'h0000000000000280;
assign   tb_i_plaintext[213]                  =   tb_i_plaintext[212];
assign   tb_o_valid[213]                      =   1'b0;
assign   tb_o_sop[213]                        =   1'b0;
assign   tb_o_ciphertext[213]                 =   tb_o_ciphertext[212];
assign   tb_o_tag_ready[213]                  =   1'b0;
assign   tb_o_tag[213]                        =   tb_o_tag[212];

// CLK no. 214/1240
// *************************************************
assign   tb_i_valid[214]                      =   1'b0;
assign   tb_i_reset[214]                      =   1'b0;
assign   tb_i_sop[214]                        =   1'b0;
assign   tb_i_key_update[214]                 =   1'b0;
assign   tb_i_key[214]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[214]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[214]               =   1'b0;
assign   tb_i_rf_static_encrypt[214]          =   1'b1;
assign   tb_i_clear_fault_flags[214]          =   1'b0;
assign   tb_i_rf_static_aad_length[214]       =   64'h0000000000000100;
assign   tb_i_aad[214]                        =   tb_i_aad[213];
assign   tb_i_rf_static_plaintext_length[214] =   64'h0000000000000280;
assign   tb_i_plaintext[214]                  =   tb_i_plaintext[213];
assign   tb_o_valid[214]                      =   1'b0;
assign   tb_o_sop[214]                        =   1'b0;
assign   tb_o_ciphertext[214]                 =   tb_o_ciphertext[213];
assign   tb_o_tag_ready[214]                  =   1'b0;
assign   tb_o_tag[214]                        =   tb_o_tag[213];

// CLK no. 215/1240
// *************************************************
assign   tb_i_valid[215]                      =   1'b0;
assign   tb_i_reset[215]                      =   1'b0;
assign   tb_i_sop[215]                        =   1'b0;
assign   tb_i_key_update[215]                 =   1'b0;
assign   tb_i_key[215]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[215]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[215]               =   1'b0;
assign   tb_i_rf_static_encrypt[215]          =   1'b1;
assign   tb_i_clear_fault_flags[215]          =   1'b0;
assign   tb_i_rf_static_aad_length[215]       =   64'h0000000000000100;
assign   tb_i_aad[215]                        =   tb_i_aad[214];
assign   tb_i_rf_static_plaintext_length[215] =   64'h0000000000000280;
assign   tb_i_plaintext[215]                  =   tb_i_plaintext[214];
assign   tb_o_valid[215]                      =   1'b0;
assign   tb_o_sop[215]                        =   1'b0;
assign   tb_o_ciphertext[215]                 =   tb_o_ciphertext[214];
assign   tb_o_tag_ready[215]                  =   1'b0;
assign   tb_o_tag[215]                        =   tb_o_tag[214];

// CLK no. 216/1240
// *************************************************
assign   tb_i_valid[216]                      =   1'b0;
assign   tb_i_reset[216]                      =   1'b0;
assign   tb_i_sop[216]                        =   1'b0;
assign   tb_i_key_update[216]                 =   1'b0;
assign   tb_i_key[216]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[216]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[216]               =   1'b0;
assign   tb_i_rf_static_encrypt[216]          =   1'b1;
assign   tb_i_clear_fault_flags[216]          =   1'b0;
assign   tb_i_rf_static_aad_length[216]       =   64'h0000000000000100;
assign   tb_i_aad[216]                        =   tb_i_aad[215];
assign   tb_i_rf_static_plaintext_length[216] =   64'h0000000000000280;
assign   tb_i_plaintext[216]                  =   tb_i_plaintext[215];
assign   tb_o_valid[216]                      =   1'b0;
assign   tb_o_sop[216]                        =   1'b0;
assign   tb_o_ciphertext[216]                 =   tb_o_ciphertext[215];
assign   tb_o_tag_ready[216]                  =   1'b0;
assign   tb_o_tag[216]                        =   tb_o_tag[215];

// CLK no. 217/1240
// *************************************************
assign   tb_i_valid[217]                      =   1'b0;
assign   tb_i_reset[217]                      =   1'b0;
assign   tb_i_sop[217]                        =   1'b0;
assign   tb_i_key_update[217]                 =   1'b0;
assign   tb_i_key[217]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[217]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[217]               =   1'b0;
assign   tb_i_rf_static_encrypt[217]          =   1'b1;
assign   tb_i_clear_fault_flags[217]          =   1'b0;
assign   tb_i_rf_static_aad_length[217]       =   64'h0000000000000100;
assign   tb_i_aad[217]                        =   tb_i_aad[216];
assign   tb_i_rf_static_plaintext_length[217] =   64'h0000000000000280;
assign   tb_i_plaintext[217]                  =   tb_i_plaintext[216];
assign   tb_o_valid[217]                      =   1'b0;
assign   tb_o_sop[217]                        =   1'b0;
assign   tb_o_ciphertext[217]                 =   tb_o_ciphertext[216];
assign   tb_o_tag_ready[217]                  =   1'b0;
assign   tb_o_tag[217]                        =   tb_o_tag[216];

// CLK no. 218/1240
// *************************************************
assign   tb_i_valid[218]                      =   1'b0;
assign   tb_i_reset[218]                      =   1'b0;
assign   tb_i_sop[218]                        =   1'b0;
assign   tb_i_key_update[218]                 =   1'b0;
assign   tb_i_key[218]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[218]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[218]               =   1'b0;
assign   tb_i_rf_static_encrypt[218]          =   1'b1;
assign   tb_i_clear_fault_flags[218]          =   1'b0;
assign   tb_i_rf_static_aad_length[218]       =   64'h0000000000000100;
assign   tb_i_aad[218]                        =   tb_i_aad[217];
assign   tb_i_rf_static_plaintext_length[218] =   64'h0000000000000280;
assign   tb_i_plaintext[218]                  =   tb_i_plaintext[217];
assign   tb_o_valid[218]                      =   1'b0;
assign   tb_o_sop[218]                        =   1'b0;
assign   tb_o_ciphertext[218]                 =   tb_o_ciphertext[217];
assign   tb_o_tag_ready[218]                  =   1'b0;
assign   tb_o_tag[218]                        =   tb_o_tag[217];

// CLK no. 219/1240
// *************************************************
assign   tb_i_valid[219]                      =   1'b0;
assign   tb_i_reset[219]                      =   1'b0;
assign   tb_i_sop[219]                        =   1'b0;
assign   tb_i_key_update[219]                 =   1'b0;
assign   tb_i_key[219]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[219]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[219]               =   1'b0;
assign   tb_i_rf_static_encrypt[219]          =   1'b1;
assign   tb_i_clear_fault_flags[219]          =   1'b0;
assign   tb_i_rf_static_aad_length[219]       =   64'h0000000000000100;
assign   tb_i_aad[219]                        =   tb_i_aad[218];
assign   tb_i_rf_static_plaintext_length[219] =   64'h0000000000000280;
assign   tb_i_plaintext[219]                  =   tb_i_plaintext[218];
assign   tb_o_valid[219]                      =   1'b0;
assign   tb_o_sop[219]                        =   1'b0;
assign   tb_o_ciphertext[219]                 =   tb_o_ciphertext[218];
assign   tb_o_tag_ready[219]                  =   1'b0;
assign   tb_o_tag[219]                        =   tb_o_tag[218];

// CLK no. 220/1240
// *************************************************
assign   tb_i_valid[220]                      =   1'b0;
assign   tb_i_reset[220]                      =   1'b0;
assign   tb_i_sop[220]                        =   1'b0;
assign   tb_i_key_update[220]                 =   1'b0;
assign   tb_i_key[220]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[220]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[220]               =   1'b0;
assign   tb_i_rf_static_encrypt[220]          =   1'b1;
assign   tb_i_clear_fault_flags[220]          =   1'b0;
assign   tb_i_rf_static_aad_length[220]       =   64'h0000000000000100;
assign   tb_i_aad[220]                        =   tb_i_aad[219];
assign   tb_i_rf_static_plaintext_length[220] =   64'h0000000000000280;
assign   tb_i_plaintext[220]                  =   tb_i_plaintext[219];
assign   tb_o_valid[220]                      =   1'b0;
assign   tb_o_sop[220]                        =   1'b0;
assign   tb_o_ciphertext[220]                 =   tb_o_ciphertext[219];
assign   tb_o_tag_ready[220]                  =   1'b0;
assign   tb_o_tag[220]                        =   tb_o_tag[219];

// CLK no. 221/1240
// *************************************************
assign   tb_i_valid[221]                      =   1'b0;
assign   tb_i_reset[221]                      =   1'b0;
assign   tb_i_sop[221]                        =   1'b0;
assign   tb_i_key_update[221]                 =   1'b0;
assign   tb_i_key[221]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[221]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[221]               =   1'b0;
assign   tb_i_rf_static_encrypt[221]          =   1'b1;
assign   tb_i_clear_fault_flags[221]          =   1'b0;
assign   tb_i_rf_static_aad_length[221]       =   64'h0000000000000100;
assign   tb_i_aad[221]                        =   tb_i_aad[220];
assign   tb_i_rf_static_plaintext_length[221] =   64'h0000000000000280;
assign   tb_i_plaintext[221]                  =   tb_i_plaintext[220];
assign   tb_o_valid[221]                      =   1'b0;
assign   tb_o_sop[221]                        =   1'b0;
assign   tb_o_ciphertext[221]                 =   tb_o_ciphertext[220];
assign   tb_o_tag_ready[221]                  =   1'b0;
assign   tb_o_tag[221]                        =   tb_o_tag[220];

// CLK no. 222/1240
// *************************************************
assign   tb_i_valid[222]                      =   1'b0;
assign   tb_i_reset[222]                      =   1'b0;
assign   tb_i_sop[222]                        =   1'b0;
assign   tb_i_key_update[222]                 =   1'b0;
assign   tb_i_key[222]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[222]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[222]               =   1'b0;
assign   tb_i_rf_static_encrypt[222]          =   1'b1;
assign   tb_i_clear_fault_flags[222]          =   1'b0;
assign   tb_i_rf_static_aad_length[222]       =   64'h0000000000000100;
assign   tb_i_aad[222]                        =   tb_i_aad[221];
assign   tb_i_rf_static_plaintext_length[222] =   64'h0000000000000280;
assign   tb_i_plaintext[222]                  =   tb_i_plaintext[221];
assign   tb_o_valid[222]                      =   1'b0;
assign   tb_o_sop[222]                        =   1'b0;
assign   tb_o_ciphertext[222]                 =   tb_o_ciphertext[221];
assign   tb_o_tag_ready[222]                  =   1'b0;
assign   tb_o_tag[222]                        =   tb_o_tag[221];

// CLK no. 223/1240
// *************************************************
assign   tb_i_valid[223]                      =   1'b0;
assign   tb_i_reset[223]                      =   1'b0;
assign   tb_i_sop[223]                        =   1'b0;
assign   tb_i_key_update[223]                 =   1'b0;
assign   tb_i_key[223]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[223]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[223]               =   1'b0;
assign   tb_i_rf_static_encrypt[223]          =   1'b1;
assign   tb_i_clear_fault_flags[223]          =   1'b0;
assign   tb_i_rf_static_aad_length[223]       =   64'h0000000000000100;
assign   tb_i_aad[223]                        =   tb_i_aad[222];
assign   tb_i_rf_static_plaintext_length[223] =   64'h0000000000000280;
assign   tb_i_plaintext[223]                  =   tb_i_plaintext[222];
assign   tb_o_valid[223]                      =   1'b0;
assign   tb_o_sop[223]                        =   1'b0;
assign   tb_o_ciphertext[223]                 =   tb_o_ciphertext[222];
assign   tb_o_tag_ready[223]                  =   1'b0;
assign   tb_o_tag[223]                        =   tb_o_tag[222];

// CLK no. 224/1240
// *************************************************
assign   tb_i_valid[224]                      =   1'b0;
assign   tb_i_reset[224]                      =   1'b0;
assign   tb_i_sop[224]                        =   1'b0;
assign   tb_i_key_update[224]                 =   1'b0;
assign   tb_i_key[224]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[224]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[224]               =   1'b0;
assign   tb_i_rf_static_encrypt[224]          =   1'b1;
assign   tb_i_clear_fault_flags[224]          =   1'b0;
assign   tb_i_rf_static_aad_length[224]       =   64'h0000000000000100;
assign   tb_i_aad[224]                        =   tb_i_aad[223];
assign   tb_i_rf_static_plaintext_length[224] =   64'h0000000000000280;
assign   tb_i_plaintext[224]                  =   tb_i_plaintext[223];
assign   tb_o_valid[224]                      =   1'b1;
assign   tb_o_sop[224]                        =   1'b1;
assign   tb_o_ciphertext[224]                 =   256'h1e7e27992f696adb626a887b76557180f08f2c2773f193d596d0eb05ef913b09;
assign   tb_o_tag_ready[224]                  =   1'b0;
assign   tb_o_tag[224]                        =   tb_o_tag[223];

// CLK no. 225/1240
// *************************************************
assign   tb_i_valid[225]                      =   1'b0;
assign   tb_i_reset[225]                      =   1'b0;
assign   tb_i_sop[225]                        =   1'b0;
assign   tb_i_key_update[225]                 =   1'b0;
assign   tb_i_key[225]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[225]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[225]               =   1'b0;
assign   tb_i_rf_static_encrypt[225]          =   1'b1;
assign   tb_i_clear_fault_flags[225]          =   1'b0;
assign   tb_i_rf_static_aad_length[225]       =   64'h0000000000000100;
assign   tb_i_aad[225]                        =   tb_i_aad[224];
assign   tb_i_rf_static_plaintext_length[225] =   64'h0000000000000280;
assign   tb_i_plaintext[225]                  =   tb_i_plaintext[224];
assign   tb_o_valid[225]                      =   1'b1;
assign   tb_o_sop[225]                        =   1'b0;
assign   tb_o_ciphertext[225]                 =   256'h1a34d482d4c8ac5961837e8562aacc4bba5ae504fe2b937eb52083ad5b36b20e;
assign   tb_o_tag_ready[225]                  =   1'b0;
assign   tb_o_tag[225]                        =   tb_o_tag[224];

// CLK no. 226/1240
// *************************************************
assign   tb_i_valid[226]                      =   1'b0;
assign   tb_i_reset[226]                      =   1'b0;
assign   tb_i_sop[226]                        =   1'b0;
assign   tb_i_key_update[226]                 =   1'b0;
assign   tb_i_key[226]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[226]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[226]               =   1'b0;
assign   tb_i_rf_static_encrypt[226]          =   1'b1;
assign   tb_i_clear_fault_flags[226]          =   1'b0;
assign   tb_i_rf_static_aad_length[226]       =   64'h0000000000000100;
assign   tb_i_aad[226]                        =   tb_i_aad[225];
assign   tb_i_rf_static_plaintext_length[226] =   64'h0000000000000280;
assign   tb_i_plaintext[226]                  =   tb_i_plaintext[225];
assign   tb_o_valid[226]                      =   1'b1;
assign   tb_o_sop[226]                        =   1'b0;
assign   tb_o_ciphertext[226]                 =   256'h7613de30d1e40487865411952a1742a4;
assign   tb_o_tag_ready[226]                  =   1'b0;
assign   tb_o_tag[226]                        =   tb_o_tag[225];

// CLK no. 227/1240
// *************************************************
assign   tb_i_valid[227]                      =   1'b0;
assign   tb_i_reset[227]                      =   1'b0;
assign   tb_i_sop[227]                        =   1'b0;
assign   tb_i_key_update[227]                 =   1'b0;
assign   tb_i_key[227]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[227]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[227]               =   1'b0;
assign   tb_i_rf_static_encrypt[227]          =   1'b1;
assign   tb_i_clear_fault_flags[227]          =   1'b0;
assign   tb_i_rf_static_aad_length[227]       =   64'h0000000000000100;
assign   tb_i_aad[227]                        =   tb_i_aad[226];
assign   tb_i_rf_static_plaintext_length[227] =   64'h0000000000000280;
assign   tb_i_plaintext[227]                  =   tb_i_plaintext[226];
assign   tb_o_valid[227]                      =   1'b0;
assign   tb_o_sop[227]                        =   1'b0;
assign   tb_o_ciphertext[227]                 =   tb_o_ciphertext[226];
assign   tb_o_tag_ready[227]                  =   1'b0;
assign   tb_o_tag[227]                        =   tb_o_tag[226];

// CLK no. 228/1240
// *************************************************
assign   tb_i_valid[228]                      =   1'b0;
assign   tb_i_reset[228]                      =   1'b0;
assign   tb_i_sop[228]                        =   1'b0;
assign   tb_i_key_update[228]                 =   1'b0;
assign   tb_i_key[228]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[228]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[228]               =   1'b0;
assign   tb_i_rf_static_encrypt[228]          =   1'b1;
assign   tb_i_clear_fault_flags[228]          =   1'b0;
assign   tb_i_rf_static_aad_length[228]       =   64'h0000000000000100;
assign   tb_i_aad[228]                        =   tb_i_aad[227];
assign   tb_i_rf_static_plaintext_length[228] =   64'h0000000000000280;
assign   tb_i_plaintext[228]                  =   tb_i_plaintext[227];
assign   tb_o_valid[228]                      =   1'b0;
assign   tb_o_sop[228]                        =   1'b0;
assign   tb_o_ciphertext[228]                 =   tb_o_ciphertext[227];
assign   tb_o_tag_ready[228]                  =   1'b0;
assign   tb_o_tag[228]                        =   tb_o_tag[227];

// CLK no. 229/1240
// *************************************************
assign   tb_i_valid[229]                      =   1'b0;
assign   tb_i_reset[229]                      =   1'b0;
assign   tb_i_sop[229]                        =   1'b0;
assign   tb_i_key_update[229]                 =   1'b0;
assign   tb_i_key[229]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[229]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[229]               =   1'b0;
assign   tb_i_rf_static_encrypt[229]          =   1'b1;
assign   tb_i_clear_fault_flags[229]          =   1'b0;
assign   tb_i_rf_static_aad_length[229]       =   64'h0000000000000100;
assign   tb_i_aad[229]                        =   tb_i_aad[228];
assign   tb_i_rf_static_plaintext_length[229] =   64'h0000000000000280;
assign   tb_i_plaintext[229]                  =   tb_i_plaintext[228];
assign   tb_o_valid[229]                      =   1'b0;
assign   tb_o_sop[229]                        =   1'b0;
assign   tb_o_ciphertext[229]                 =   tb_o_ciphertext[228];
assign   tb_o_tag_ready[229]                  =   1'b0;
assign   tb_o_tag[229]                        =   tb_o_tag[228];

// CLK no. 230/1240
// *************************************************
assign   tb_i_valid[230]                      =   1'b0;
assign   tb_i_reset[230]                      =   1'b0;
assign   tb_i_sop[230]                        =   1'b0;
assign   tb_i_key_update[230]                 =   1'b0;
assign   tb_i_key[230]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[230]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[230]               =   1'b0;
assign   tb_i_rf_static_encrypt[230]          =   1'b1;
assign   tb_i_clear_fault_flags[230]          =   1'b0;
assign   tb_i_rf_static_aad_length[230]       =   64'h0000000000000100;
assign   tb_i_aad[230]                        =   tb_i_aad[229];
assign   tb_i_rf_static_plaintext_length[230] =   64'h0000000000000280;
assign   tb_i_plaintext[230]                  =   tb_i_plaintext[229];
assign   tb_o_valid[230]                      =   1'b0;
assign   tb_o_sop[230]                        =   1'b0;
assign   tb_o_ciphertext[230]                 =   tb_o_ciphertext[229];
assign   tb_o_tag_ready[230]                  =   1'b0;
assign   tb_o_tag[230]                        =   tb_o_tag[229];

// CLK no. 231/1240
// *************************************************
assign   tb_i_valid[231]                      =   1'b0;
assign   tb_i_reset[231]                      =   1'b0;
assign   tb_i_sop[231]                        =   1'b0;
assign   tb_i_key_update[231]                 =   1'b0;
assign   tb_i_key[231]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[231]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[231]               =   1'b0;
assign   tb_i_rf_static_encrypt[231]          =   1'b1;
assign   tb_i_clear_fault_flags[231]          =   1'b0;
assign   tb_i_rf_static_aad_length[231]       =   64'h0000000000000100;
assign   tb_i_aad[231]                        =   tb_i_aad[230];
assign   tb_i_rf_static_plaintext_length[231] =   64'h0000000000000280;
assign   tb_i_plaintext[231]                  =   tb_i_plaintext[230];
assign   tb_o_valid[231]                      =   1'b0;
assign   tb_o_sop[231]                        =   1'b0;
assign   tb_o_ciphertext[231]                 =   tb_o_ciphertext[230];
assign   tb_o_tag_ready[231]                  =   1'b0;
assign   tb_o_tag[231]                        =   tb_o_tag[230];

// CLK no. 232/1240
// *************************************************
assign   tb_i_valid[232]                      =   1'b0;
assign   tb_i_reset[232]                      =   1'b0;
assign   tb_i_sop[232]                        =   1'b0;
assign   tb_i_key_update[232]                 =   1'b0;
assign   tb_i_key[232]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[232]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[232]               =   1'b0;
assign   tb_i_rf_static_encrypt[232]          =   1'b1;
assign   tb_i_clear_fault_flags[232]          =   1'b0;
assign   tb_i_rf_static_aad_length[232]       =   64'h0000000000000100;
assign   tb_i_aad[232]                        =   tb_i_aad[231];
assign   tb_i_rf_static_plaintext_length[232] =   64'h0000000000000280;
assign   tb_i_plaintext[232]                  =   tb_i_plaintext[231];
assign   tb_o_valid[232]                      =   1'b0;
assign   tb_o_sop[232]                        =   1'b0;
assign   tb_o_ciphertext[232]                 =   tb_o_ciphertext[231];
assign   tb_o_tag_ready[232]                  =   1'b0;
assign   tb_o_tag[232]                        =   tb_o_tag[231];

// CLK no. 233/1240
// *************************************************
assign   tb_i_valid[233]                      =   1'b0;
assign   tb_i_reset[233]                      =   1'b0;
assign   tb_i_sop[233]                        =   1'b0;
assign   tb_i_key_update[233]                 =   1'b0;
assign   tb_i_key[233]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[233]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[233]               =   1'b0;
assign   tb_i_rf_static_encrypt[233]          =   1'b1;
assign   tb_i_clear_fault_flags[233]          =   1'b0;
assign   tb_i_rf_static_aad_length[233]       =   64'h0000000000000100;
assign   tb_i_aad[233]                        =   tb_i_aad[232];
assign   tb_i_rf_static_plaintext_length[233] =   64'h0000000000000280;
assign   tb_i_plaintext[233]                  =   tb_i_plaintext[232];
assign   tb_o_valid[233]                      =   1'b0;
assign   tb_o_sop[233]                        =   1'b0;
assign   tb_o_ciphertext[233]                 =   tb_o_ciphertext[232];
assign   tb_o_tag_ready[233]                  =   1'b0;
assign   tb_o_tag[233]                        =   tb_o_tag[232];

// CLK no. 234/1240
// *************************************************
assign   tb_i_valid[234]                      =   1'b0;
assign   tb_i_reset[234]                      =   1'b0;
assign   tb_i_sop[234]                        =   1'b0;
assign   tb_i_key_update[234]                 =   1'b0;
assign   tb_i_key[234]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[234]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[234]               =   1'b0;
assign   tb_i_rf_static_encrypt[234]          =   1'b1;
assign   tb_i_clear_fault_flags[234]          =   1'b0;
assign   tb_i_rf_static_aad_length[234]       =   64'h0000000000000100;
assign   tb_i_aad[234]                        =   tb_i_aad[233];
assign   tb_i_rf_static_plaintext_length[234] =   64'h0000000000000280;
assign   tb_i_plaintext[234]                  =   tb_i_plaintext[233];
assign   tb_o_valid[234]                      =   1'b0;
assign   tb_o_sop[234]                        =   1'b0;
assign   tb_o_ciphertext[234]                 =   tb_o_ciphertext[233];
assign   tb_o_tag_ready[234]                  =   1'b1;
assign   tb_o_tag[234]                        =   128'h3b52ba731b51aa92f8939014a047fab9;

// CLK no. 235/1240
// *************************************************
assign   tb_i_valid[235]                      =   1'b0;
assign   tb_i_reset[235]                      =   1'b0;
assign   tb_i_sop[235]                        =   1'b0;
assign   tb_i_key_update[235]                 =   1'b0;
assign   tb_i_key[235]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[235]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[235]               =   1'b0;
assign   tb_i_rf_static_encrypt[235]          =   1'b1;
assign   tb_i_clear_fault_flags[235]          =   1'b0;
assign   tb_i_rf_static_aad_length[235]       =   64'h0000000000000100;
assign   tb_i_aad[235]                        =   tb_i_aad[234];
assign   tb_i_rf_static_plaintext_length[235] =   64'h0000000000000280;
assign   tb_i_plaintext[235]                  =   tb_i_plaintext[234];
assign   tb_o_valid[235]                      =   1'b0;
assign   tb_o_sop[235]                        =   1'b0;
assign   tb_o_ciphertext[235]                 =   tb_o_ciphertext[234];
assign   tb_o_tag_ready[235]                  =   1'b0;
assign   tb_o_tag[235]                        =   tb_o_tag[234];

// CLK no. 236/1240
// *************************************************
assign   tb_i_valid[236]                      =   1'b0;
assign   tb_i_reset[236]                      =   1'b0;
assign   tb_i_sop[236]                        =   1'b0;
assign   tb_i_key_update[236]                 =   1'b0;
assign   tb_i_key[236]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[236]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[236]               =   1'b0;
assign   tb_i_rf_static_encrypt[236]          =   1'b1;
assign   tb_i_clear_fault_flags[236]          =   1'b0;
assign   tb_i_rf_static_aad_length[236]       =   64'h0000000000000100;
assign   tb_i_aad[236]                        =   tb_i_aad[235];
assign   tb_i_rf_static_plaintext_length[236] =   64'h0000000000000280;
assign   tb_i_plaintext[236]                  =   tb_i_plaintext[235];
assign   tb_o_valid[236]                      =   1'b0;
assign   tb_o_sop[236]                        =   1'b0;
assign   tb_o_ciphertext[236]                 =   tb_o_ciphertext[235];
assign   tb_o_tag_ready[236]                  =   1'b0;
assign   tb_o_tag[236]                        =   tb_o_tag[235];

// CLK no. 237/1240
// *************************************************
assign   tb_i_valid[237]                      =   1'b0;
assign   tb_i_reset[237]                      =   1'b0;
assign   tb_i_sop[237]                        =   1'b1;
assign   tb_i_key_update[237]                 =   1'b0;
assign   tb_i_key[237]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[237]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[237]               =   1'b0;
assign   tb_i_rf_static_encrypt[237]          =   1'b1;
assign   tb_i_clear_fault_flags[237]          =   1'b0;
assign   tb_i_rf_static_aad_length[237]       =   64'h0000000000000100;
assign   tb_i_aad[237]                        =   tb_i_aad[236];
assign   tb_i_rf_static_plaintext_length[237] =   64'h0000000000000280;
assign   tb_i_plaintext[237]                  =   tb_i_plaintext[236];
assign   tb_o_valid[237]                      =   1'b0;
assign   tb_o_sop[237]                        =   1'b0;
assign   tb_o_ciphertext[237]                 =   tb_o_ciphertext[236];
assign   tb_o_tag_ready[237]                  =   1'b0;
assign   tb_o_tag[237]                        =   tb_o_tag[236];

// CLK no. 238/1240
// *************************************************
assign   tb_i_valid[238]                      =   1'b1;
assign   tb_i_reset[238]                      =   1'b0;
assign   tb_i_sop[238]                        =   1'b0;
assign   tb_i_key_update[238]                 =   1'b0;
assign   tb_i_key[238]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[238]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[238]               =   1'b0;
assign   tb_i_rf_static_encrypt[238]          =   1'b1;
assign   tb_i_clear_fault_flags[238]          =   1'b0;
assign   tb_i_rf_static_aad_length[238]       =   64'h0000000000000100;
assign   tb_i_aad[238]                        =   256'h366cd9ed8f74a477b61c41296282d756827e64811b319cc1cb9b0a494bec4a15;
assign   tb_i_rf_static_plaintext_length[238] =   64'h0000000000000280;
assign   tb_i_plaintext[238]                  =   tb_i_plaintext[237];
assign   tb_o_valid[238]                      =   1'b0;
assign   tb_o_sop[238]                        =   1'b0;
assign   tb_o_ciphertext[238]                 =   tb_o_ciphertext[237];
assign   tb_o_tag_ready[238]                  =   1'b0;
assign   tb_o_tag[238]                        =   tb_o_tag[237];

// CLK no. 239/1240
// *************************************************
assign   tb_i_valid[239]                      =   1'b1;
assign   tb_i_reset[239]                      =   1'b0;
assign   tb_i_sop[239]                        =   1'b0;
assign   tb_i_key_update[239]                 =   1'b0;
assign   tb_i_key[239]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[239]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[239]               =   1'b0;
assign   tb_i_rf_static_encrypt[239]          =   1'b1;
assign   tb_i_clear_fault_flags[239]          =   1'b0;
assign   tb_i_rf_static_aad_length[239]       =   64'h0000000000000100;
assign   tb_i_aad[239]                        =   tb_i_aad[238];
assign   tb_i_rf_static_plaintext_length[239] =   64'h0000000000000280;
assign   tb_i_plaintext[239]                  =   256'h6564939754d1d738def6d459de6479c16a461a9bd961680f19bd94a46c4ee246;
assign   tb_o_valid[239]                      =   1'b0;
assign   tb_o_sop[239]                        =   1'b0;
assign   tb_o_ciphertext[239]                 =   tb_o_ciphertext[238];
assign   tb_o_tag_ready[239]                  =   1'b0;
assign   tb_o_tag[239]                        =   tb_o_tag[238];

// CLK no. 240/1240
// *************************************************
assign   tb_i_valid[240]                      =   1'b1;
assign   tb_i_reset[240]                      =   1'b0;
assign   tb_i_sop[240]                        =   1'b0;
assign   tb_i_key_update[240]                 =   1'b0;
assign   tb_i_key[240]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[240]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[240]               =   1'b0;
assign   tb_i_rf_static_encrypt[240]          =   1'b1;
assign   tb_i_clear_fault_flags[240]          =   1'b0;
assign   tb_i_rf_static_aad_length[240]       =   64'h0000000000000100;
assign   tb_i_aad[240]                        =   tb_i_aad[239];
assign   tb_i_rf_static_plaintext_length[240] =   64'h0000000000000280;
assign   tb_i_plaintext[240]                  =   256'hb8b5e9686e8275170678cc8550fef8c6852c487f4f9e2cb8667ae4b847f864bf;
assign   tb_o_valid[240]                      =   1'b0;
assign   tb_o_sop[240]                        =   1'b0;
assign   tb_o_ciphertext[240]                 =   tb_o_ciphertext[239];
assign   tb_o_tag_ready[240]                  =   1'b0;
assign   tb_o_tag[240]                        =   tb_o_tag[239];

// CLK no. 241/1240
// *************************************************
assign   tb_i_valid[241]                      =   1'b1;
assign   tb_i_reset[241]                      =   1'b0;
assign   tb_i_sop[241]                        =   1'b0;
assign   tb_i_key_update[241]                 =   1'b0;
assign   tb_i_key[241]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[241]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[241]               =   1'b0;
assign   tb_i_rf_static_encrypt[241]          =   1'b1;
assign   tb_i_clear_fault_flags[241]          =   1'b0;
assign   tb_i_rf_static_aad_length[241]       =   64'h0000000000000100;
assign   tb_i_aad[241]                        =   tb_i_aad[240];
assign   tb_i_rf_static_plaintext_length[241] =   64'h0000000000000280;
assign   tb_i_plaintext[241]                  =   256'hbcd4183e647b475b380b9a14925fa35a;
assign   tb_o_valid[241]                      =   1'b0;
assign   tb_o_sop[241]                        =   1'b0;
assign   tb_o_ciphertext[241]                 =   tb_o_ciphertext[240];
assign   tb_o_tag_ready[241]                  =   1'b0;
assign   tb_o_tag[241]                        =   tb_o_tag[240];

// CLK no. 242/1240
// *************************************************
assign   tb_i_valid[242]                      =   1'b0;
assign   tb_i_reset[242]                      =   1'b0;
assign   tb_i_sop[242]                        =   1'b0;
assign   tb_i_key_update[242]                 =   1'b0;
assign   tb_i_key[242]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[242]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[242]               =   1'b0;
assign   tb_i_rf_static_encrypt[242]          =   1'b1;
assign   tb_i_clear_fault_flags[242]          =   1'b0;
assign   tb_i_rf_static_aad_length[242]       =   64'h0000000000000100;
assign   tb_i_aad[242]                        =   tb_i_aad[241];
assign   tb_i_rf_static_plaintext_length[242] =   64'h0000000000000280;
assign   tb_i_plaintext[242]                  =   tb_i_plaintext[241];
assign   tb_o_valid[242]                      =   1'b0;
assign   tb_o_sop[242]                        =   1'b0;
assign   tb_o_ciphertext[242]                 =   tb_o_ciphertext[241];
assign   tb_o_tag_ready[242]                  =   1'b0;
assign   tb_o_tag[242]                        =   tb_o_tag[241];

// CLK no. 243/1240
// *************************************************
assign   tb_i_valid[243]                      =   1'b0;
assign   tb_i_reset[243]                      =   1'b0;
assign   tb_i_sop[243]                        =   1'b0;
assign   tb_i_key_update[243]                 =   1'b0;
assign   tb_i_key[243]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[243]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[243]               =   1'b0;
assign   tb_i_rf_static_encrypt[243]          =   1'b1;
assign   tb_i_clear_fault_flags[243]          =   1'b0;
assign   tb_i_rf_static_aad_length[243]       =   64'h0000000000000100;
assign   tb_i_aad[243]                        =   tb_i_aad[242];
assign   tb_i_rf_static_plaintext_length[243] =   64'h0000000000000280;
assign   tb_i_plaintext[243]                  =   tb_i_plaintext[242];
assign   tb_o_valid[243]                      =   1'b0;
assign   tb_o_sop[243]                        =   1'b0;
assign   tb_o_ciphertext[243]                 =   tb_o_ciphertext[242];
assign   tb_o_tag_ready[243]                  =   1'b0;
assign   tb_o_tag[243]                        =   tb_o_tag[242];

// CLK no. 244/1240
// *************************************************
assign   tb_i_valid[244]                      =   1'b0;
assign   tb_i_reset[244]                      =   1'b0;
assign   tb_i_sop[244]                        =   1'b0;
assign   tb_i_key_update[244]                 =   1'b0;
assign   tb_i_key[244]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[244]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[244]               =   1'b0;
assign   tb_i_rf_static_encrypt[244]          =   1'b1;
assign   tb_i_clear_fault_flags[244]          =   1'b0;
assign   tb_i_rf_static_aad_length[244]       =   64'h0000000000000100;
assign   tb_i_aad[244]                        =   tb_i_aad[243];
assign   tb_i_rf_static_plaintext_length[244] =   64'h0000000000000280;
assign   tb_i_plaintext[244]                  =   tb_i_plaintext[243];
assign   tb_o_valid[244]                      =   1'b0;
assign   tb_o_sop[244]                        =   1'b0;
assign   tb_o_ciphertext[244]                 =   tb_o_ciphertext[243];
assign   tb_o_tag_ready[244]                  =   1'b0;
assign   tb_o_tag[244]                        =   tb_o_tag[243];

// CLK no. 245/1240
// *************************************************
assign   tb_i_valid[245]                      =   1'b0;
assign   tb_i_reset[245]                      =   1'b0;
assign   tb_i_sop[245]                        =   1'b0;
assign   tb_i_key_update[245]                 =   1'b0;
assign   tb_i_key[245]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[245]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[245]               =   1'b0;
assign   tb_i_rf_static_encrypt[245]          =   1'b1;
assign   tb_i_clear_fault_flags[245]          =   1'b0;
assign   tb_i_rf_static_aad_length[245]       =   64'h0000000000000100;
assign   tb_i_aad[245]                        =   tb_i_aad[244];
assign   tb_i_rf_static_plaintext_length[245] =   64'h0000000000000280;
assign   tb_i_plaintext[245]                  =   tb_i_plaintext[244];
assign   tb_o_valid[245]                      =   1'b0;
assign   tb_o_sop[245]                        =   1'b0;
assign   tb_o_ciphertext[245]                 =   tb_o_ciphertext[244];
assign   tb_o_tag_ready[245]                  =   1'b0;
assign   tb_o_tag[245]                        =   tb_o_tag[244];

// CLK no. 246/1240
// *************************************************
assign   tb_i_valid[246]                      =   1'b0;
assign   tb_i_reset[246]                      =   1'b0;
assign   tb_i_sop[246]                        =   1'b0;
assign   tb_i_key_update[246]                 =   1'b0;
assign   tb_i_key[246]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[246]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[246]               =   1'b0;
assign   tb_i_rf_static_encrypt[246]          =   1'b1;
assign   tb_i_clear_fault_flags[246]          =   1'b0;
assign   tb_i_rf_static_aad_length[246]       =   64'h0000000000000100;
assign   tb_i_aad[246]                        =   tb_i_aad[245];
assign   tb_i_rf_static_plaintext_length[246] =   64'h0000000000000280;
assign   tb_i_plaintext[246]                  =   tb_i_plaintext[245];
assign   tb_o_valid[246]                      =   1'b0;
assign   tb_o_sop[246]                        =   1'b0;
assign   tb_o_ciphertext[246]                 =   tb_o_ciphertext[245];
assign   tb_o_tag_ready[246]                  =   1'b0;
assign   tb_o_tag[246]                        =   tb_o_tag[245];

// CLK no. 247/1240
// *************************************************
assign   tb_i_valid[247]                      =   1'b0;
assign   tb_i_reset[247]                      =   1'b0;
assign   tb_i_sop[247]                        =   1'b0;
assign   tb_i_key_update[247]                 =   1'b0;
assign   tb_i_key[247]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[247]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[247]               =   1'b0;
assign   tb_i_rf_static_encrypt[247]          =   1'b1;
assign   tb_i_clear_fault_flags[247]          =   1'b0;
assign   tb_i_rf_static_aad_length[247]       =   64'h0000000000000100;
assign   tb_i_aad[247]                        =   tb_i_aad[246];
assign   tb_i_rf_static_plaintext_length[247] =   64'h0000000000000280;
assign   tb_i_plaintext[247]                  =   tb_i_plaintext[246];
assign   tb_o_valid[247]                      =   1'b0;
assign   tb_o_sop[247]                        =   1'b0;
assign   tb_o_ciphertext[247]                 =   tb_o_ciphertext[246];
assign   tb_o_tag_ready[247]                  =   1'b0;
assign   tb_o_tag[247]                        =   tb_o_tag[246];

// CLK no. 248/1240
// *************************************************
assign   tb_i_valid[248]                      =   1'b0;
assign   tb_i_reset[248]                      =   1'b0;
assign   tb_i_sop[248]                        =   1'b0;
assign   tb_i_key_update[248]                 =   1'b0;
assign   tb_i_key[248]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[248]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[248]               =   1'b0;
assign   tb_i_rf_static_encrypt[248]          =   1'b1;
assign   tb_i_clear_fault_flags[248]          =   1'b0;
assign   tb_i_rf_static_aad_length[248]       =   64'h0000000000000100;
assign   tb_i_aad[248]                        =   tb_i_aad[247];
assign   tb_i_rf_static_plaintext_length[248] =   64'h0000000000000280;
assign   tb_i_plaintext[248]                  =   tb_i_plaintext[247];
assign   tb_o_valid[248]                      =   1'b0;
assign   tb_o_sop[248]                        =   1'b0;
assign   tb_o_ciphertext[248]                 =   tb_o_ciphertext[247];
assign   tb_o_tag_ready[248]                  =   1'b0;
assign   tb_o_tag[248]                        =   tb_o_tag[247];

// CLK no. 249/1240
// *************************************************
assign   tb_i_valid[249]                      =   1'b0;
assign   tb_i_reset[249]                      =   1'b0;
assign   tb_i_sop[249]                        =   1'b0;
assign   tb_i_key_update[249]                 =   1'b0;
assign   tb_i_key[249]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[249]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[249]               =   1'b0;
assign   tb_i_rf_static_encrypt[249]          =   1'b1;
assign   tb_i_clear_fault_flags[249]          =   1'b0;
assign   tb_i_rf_static_aad_length[249]       =   64'h0000000000000100;
assign   tb_i_aad[249]                        =   tb_i_aad[248];
assign   tb_i_rf_static_plaintext_length[249] =   64'h0000000000000280;
assign   tb_i_plaintext[249]                  =   tb_i_plaintext[248];
assign   tb_o_valid[249]                      =   1'b0;
assign   tb_o_sop[249]                        =   1'b0;
assign   tb_o_ciphertext[249]                 =   tb_o_ciphertext[248];
assign   tb_o_tag_ready[249]                  =   1'b0;
assign   tb_o_tag[249]                        =   tb_o_tag[248];

// CLK no. 250/1240
// *************************************************
assign   tb_i_valid[250]                      =   1'b0;
assign   tb_i_reset[250]                      =   1'b0;
assign   tb_i_sop[250]                        =   1'b0;
assign   tb_i_key_update[250]                 =   1'b0;
assign   tb_i_key[250]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[250]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[250]               =   1'b0;
assign   tb_i_rf_static_encrypt[250]          =   1'b1;
assign   tb_i_clear_fault_flags[250]          =   1'b0;
assign   tb_i_rf_static_aad_length[250]       =   64'h0000000000000100;
assign   tb_i_aad[250]                        =   tb_i_aad[249];
assign   tb_i_rf_static_plaintext_length[250] =   64'h0000000000000280;
assign   tb_i_plaintext[250]                  =   tb_i_plaintext[249];
assign   tb_o_valid[250]                      =   1'b0;
assign   tb_o_sop[250]                        =   1'b0;
assign   tb_o_ciphertext[250]                 =   tb_o_ciphertext[249];
assign   tb_o_tag_ready[250]                  =   1'b0;
assign   tb_o_tag[250]                        =   tb_o_tag[249];

// CLK no. 251/1240
// *************************************************
assign   tb_i_valid[251]                      =   1'b0;
assign   tb_i_reset[251]                      =   1'b0;
assign   tb_i_sop[251]                        =   1'b0;
assign   tb_i_key_update[251]                 =   1'b0;
assign   tb_i_key[251]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[251]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[251]               =   1'b0;
assign   tb_i_rf_static_encrypt[251]          =   1'b1;
assign   tb_i_clear_fault_flags[251]          =   1'b0;
assign   tb_i_rf_static_aad_length[251]       =   64'h0000000000000100;
assign   tb_i_aad[251]                        =   tb_i_aad[250];
assign   tb_i_rf_static_plaintext_length[251] =   64'h0000000000000280;
assign   tb_i_plaintext[251]                  =   tb_i_plaintext[250];
assign   tb_o_valid[251]                      =   1'b0;
assign   tb_o_sop[251]                        =   1'b0;
assign   tb_o_ciphertext[251]                 =   tb_o_ciphertext[250];
assign   tb_o_tag_ready[251]                  =   1'b0;
assign   tb_o_tag[251]                        =   tb_o_tag[250];

// CLK no. 252/1240
// *************************************************
assign   tb_i_valid[252]                      =   1'b0;
assign   tb_i_reset[252]                      =   1'b0;
assign   tb_i_sop[252]                        =   1'b0;
assign   tb_i_key_update[252]                 =   1'b0;
assign   tb_i_key[252]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[252]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[252]               =   1'b0;
assign   tb_i_rf_static_encrypt[252]          =   1'b1;
assign   tb_i_clear_fault_flags[252]          =   1'b0;
assign   tb_i_rf_static_aad_length[252]       =   64'h0000000000000100;
assign   tb_i_aad[252]                        =   tb_i_aad[251];
assign   tb_i_rf_static_plaintext_length[252] =   64'h0000000000000280;
assign   tb_i_plaintext[252]                  =   tb_i_plaintext[251];
assign   tb_o_valid[252]                      =   1'b0;
assign   tb_o_sop[252]                        =   1'b0;
assign   tb_o_ciphertext[252]                 =   tb_o_ciphertext[251];
assign   tb_o_tag_ready[252]                  =   1'b0;
assign   tb_o_tag[252]                        =   tb_o_tag[251];

// CLK no. 253/1240
// *************************************************
assign   tb_i_valid[253]                      =   1'b0;
assign   tb_i_reset[253]                      =   1'b0;
assign   tb_i_sop[253]                        =   1'b0;
assign   tb_i_key_update[253]                 =   1'b0;
assign   tb_i_key[253]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[253]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[253]               =   1'b0;
assign   tb_i_rf_static_encrypt[253]          =   1'b1;
assign   tb_i_clear_fault_flags[253]          =   1'b0;
assign   tb_i_rf_static_aad_length[253]       =   64'h0000000000000100;
assign   tb_i_aad[253]                        =   tb_i_aad[252];
assign   tb_i_rf_static_plaintext_length[253] =   64'h0000000000000280;
assign   tb_i_plaintext[253]                  =   tb_i_plaintext[252];
assign   tb_o_valid[253]                      =   1'b0;
assign   tb_o_sop[253]                        =   1'b0;
assign   tb_o_ciphertext[253]                 =   tb_o_ciphertext[252];
assign   tb_o_tag_ready[253]                  =   1'b0;
assign   tb_o_tag[253]                        =   tb_o_tag[252];

// CLK no. 254/1240
// *************************************************
assign   tb_i_valid[254]                      =   1'b0;
assign   tb_i_reset[254]                      =   1'b0;
assign   tb_i_sop[254]                        =   1'b0;
assign   tb_i_key_update[254]                 =   1'b0;
assign   tb_i_key[254]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[254]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[254]               =   1'b0;
assign   tb_i_rf_static_encrypt[254]          =   1'b1;
assign   tb_i_clear_fault_flags[254]          =   1'b0;
assign   tb_i_rf_static_aad_length[254]       =   64'h0000000000000100;
assign   tb_i_aad[254]                        =   tb_i_aad[253];
assign   tb_i_rf_static_plaintext_length[254] =   64'h0000000000000280;
assign   tb_i_plaintext[254]                  =   tb_i_plaintext[253];
assign   tb_o_valid[254]                      =   1'b0;
assign   tb_o_sop[254]                        =   1'b0;
assign   tb_o_ciphertext[254]                 =   tb_o_ciphertext[253];
assign   tb_o_tag_ready[254]                  =   1'b0;
assign   tb_o_tag[254]                        =   tb_o_tag[253];

// CLK no. 255/1240
// *************************************************
assign   tb_i_valid[255]                      =   1'b0;
assign   tb_i_reset[255]                      =   1'b0;
assign   tb_i_sop[255]                        =   1'b0;
assign   tb_i_key_update[255]                 =   1'b0;
assign   tb_i_key[255]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[255]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[255]               =   1'b0;
assign   tb_i_rf_static_encrypt[255]          =   1'b1;
assign   tb_i_clear_fault_flags[255]          =   1'b0;
assign   tb_i_rf_static_aad_length[255]       =   64'h0000000000000100;
assign   tb_i_aad[255]                        =   tb_i_aad[254];
assign   tb_i_rf_static_plaintext_length[255] =   64'h0000000000000280;
assign   tb_i_plaintext[255]                  =   tb_i_plaintext[254];
assign   tb_o_valid[255]                      =   1'b0;
assign   tb_o_sop[255]                        =   1'b0;
assign   tb_o_ciphertext[255]                 =   tb_o_ciphertext[254];
assign   tb_o_tag_ready[255]                  =   1'b0;
assign   tb_o_tag[255]                        =   tb_o_tag[254];

// CLK no. 256/1240
// *************************************************
assign   tb_i_valid[256]                      =   1'b0;
assign   tb_i_reset[256]                      =   1'b0;
assign   tb_i_sop[256]                        =   1'b0;
assign   tb_i_key_update[256]                 =   1'b0;
assign   tb_i_key[256]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[256]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[256]               =   1'b0;
assign   tb_i_rf_static_encrypt[256]          =   1'b1;
assign   tb_i_clear_fault_flags[256]          =   1'b0;
assign   tb_i_rf_static_aad_length[256]       =   64'h0000000000000100;
assign   tb_i_aad[256]                        =   tb_i_aad[255];
assign   tb_i_rf_static_plaintext_length[256] =   64'h0000000000000280;
assign   tb_i_plaintext[256]                  =   tb_i_plaintext[255];
assign   tb_o_valid[256]                      =   1'b0;
assign   tb_o_sop[256]                        =   1'b0;
assign   tb_o_ciphertext[256]                 =   tb_o_ciphertext[255];
assign   tb_o_tag_ready[256]                  =   1'b0;
assign   tb_o_tag[256]                        =   tb_o_tag[255];

// CLK no. 257/1240
// *************************************************
assign   tb_i_valid[257]                      =   1'b0;
assign   tb_i_reset[257]                      =   1'b0;
assign   tb_i_sop[257]                        =   1'b0;
assign   tb_i_key_update[257]                 =   1'b0;
assign   tb_i_key[257]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[257]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[257]               =   1'b0;
assign   tb_i_rf_static_encrypt[257]          =   1'b1;
assign   tb_i_clear_fault_flags[257]          =   1'b0;
assign   tb_i_rf_static_aad_length[257]       =   64'h0000000000000100;
assign   tb_i_aad[257]                        =   tb_i_aad[256];
assign   tb_i_rf_static_plaintext_length[257] =   64'h0000000000000280;
assign   tb_i_plaintext[257]                  =   tb_i_plaintext[256];
assign   tb_o_valid[257]                      =   1'b0;
assign   tb_o_sop[257]                        =   1'b0;
assign   tb_o_ciphertext[257]                 =   tb_o_ciphertext[256];
assign   tb_o_tag_ready[257]                  =   1'b0;
assign   tb_o_tag[257]                        =   tb_o_tag[256];

// CLK no. 258/1240
// *************************************************
assign   tb_i_valid[258]                      =   1'b0;
assign   tb_i_reset[258]                      =   1'b0;
assign   tb_i_sop[258]                        =   1'b0;
assign   tb_i_key_update[258]                 =   1'b0;
assign   tb_i_key[258]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[258]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[258]               =   1'b0;
assign   tb_i_rf_static_encrypt[258]          =   1'b1;
assign   tb_i_clear_fault_flags[258]          =   1'b0;
assign   tb_i_rf_static_aad_length[258]       =   64'h0000000000000100;
assign   tb_i_aad[258]                        =   tb_i_aad[257];
assign   tb_i_rf_static_plaintext_length[258] =   64'h0000000000000280;
assign   tb_i_plaintext[258]                  =   tb_i_plaintext[257];
assign   tb_o_valid[258]                      =   1'b0;
assign   tb_o_sop[258]                        =   1'b0;
assign   tb_o_ciphertext[258]                 =   tb_o_ciphertext[257];
assign   tb_o_tag_ready[258]                  =   1'b0;
assign   tb_o_tag[258]                        =   tb_o_tag[257];

// CLK no. 259/1240
// *************************************************
assign   tb_i_valid[259]                      =   1'b0;
assign   tb_i_reset[259]                      =   1'b0;
assign   tb_i_sop[259]                        =   1'b0;
assign   tb_i_key_update[259]                 =   1'b0;
assign   tb_i_key[259]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[259]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[259]               =   1'b0;
assign   tb_i_rf_static_encrypt[259]          =   1'b1;
assign   tb_i_clear_fault_flags[259]          =   1'b0;
assign   tb_i_rf_static_aad_length[259]       =   64'h0000000000000100;
assign   tb_i_aad[259]                        =   tb_i_aad[258];
assign   tb_i_rf_static_plaintext_length[259] =   64'h0000000000000280;
assign   tb_i_plaintext[259]                  =   tb_i_plaintext[258];
assign   tb_o_valid[259]                      =   1'b0;
assign   tb_o_sop[259]                        =   1'b0;
assign   tb_o_ciphertext[259]                 =   tb_o_ciphertext[258];
assign   tb_o_tag_ready[259]                  =   1'b0;
assign   tb_o_tag[259]                        =   tb_o_tag[258];

// CLK no. 260/1240
// *************************************************
assign   tb_i_valid[260]                      =   1'b0;
assign   tb_i_reset[260]                      =   1'b0;
assign   tb_i_sop[260]                        =   1'b0;
assign   tb_i_key_update[260]                 =   1'b0;
assign   tb_i_key[260]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[260]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[260]               =   1'b0;
assign   tb_i_rf_static_encrypt[260]          =   1'b1;
assign   tb_i_clear_fault_flags[260]          =   1'b0;
assign   tb_i_rf_static_aad_length[260]       =   64'h0000000000000100;
assign   tb_i_aad[260]                        =   tb_i_aad[259];
assign   tb_i_rf_static_plaintext_length[260] =   64'h0000000000000280;
assign   tb_i_plaintext[260]                  =   tb_i_plaintext[259];
assign   tb_o_valid[260]                      =   1'b0;
assign   tb_o_sop[260]                        =   1'b0;
assign   tb_o_ciphertext[260]                 =   tb_o_ciphertext[259];
assign   tb_o_tag_ready[260]                  =   1'b0;
assign   tb_o_tag[260]                        =   tb_o_tag[259];

// CLK no. 261/1240
// *************************************************
assign   tb_i_valid[261]                      =   1'b0;
assign   tb_i_reset[261]                      =   1'b0;
assign   tb_i_sop[261]                        =   1'b0;
assign   tb_i_key_update[261]                 =   1'b0;
assign   tb_i_key[261]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[261]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[261]               =   1'b0;
assign   tb_i_rf_static_encrypt[261]          =   1'b1;
assign   tb_i_clear_fault_flags[261]          =   1'b0;
assign   tb_i_rf_static_aad_length[261]       =   64'h0000000000000100;
assign   tb_i_aad[261]                        =   tb_i_aad[260];
assign   tb_i_rf_static_plaintext_length[261] =   64'h0000000000000280;
assign   tb_i_plaintext[261]                  =   tb_i_plaintext[260];
assign   tb_o_valid[261]                      =   1'b0;
assign   tb_o_sop[261]                        =   1'b0;
assign   tb_o_ciphertext[261]                 =   tb_o_ciphertext[260];
assign   tb_o_tag_ready[261]                  =   1'b0;
assign   tb_o_tag[261]                        =   tb_o_tag[260];

// CLK no. 262/1240
// *************************************************
assign   tb_i_valid[262]                      =   1'b0;
assign   tb_i_reset[262]                      =   1'b0;
assign   tb_i_sop[262]                        =   1'b0;
assign   tb_i_key_update[262]                 =   1'b0;
assign   tb_i_key[262]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[262]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[262]               =   1'b0;
assign   tb_i_rf_static_encrypt[262]          =   1'b1;
assign   tb_i_clear_fault_flags[262]          =   1'b0;
assign   tb_i_rf_static_aad_length[262]       =   64'h0000000000000100;
assign   tb_i_aad[262]                        =   tb_i_aad[261];
assign   tb_i_rf_static_plaintext_length[262] =   64'h0000000000000280;
assign   tb_i_plaintext[262]                  =   tb_i_plaintext[261];
assign   tb_o_valid[262]                      =   1'b0;
assign   tb_o_sop[262]                        =   1'b0;
assign   tb_o_ciphertext[262]                 =   tb_o_ciphertext[261];
assign   tb_o_tag_ready[262]                  =   1'b0;
assign   tb_o_tag[262]                        =   tb_o_tag[261];

// CLK no. 263/1240
// *************************************************
assign   tb_i_valid[263]                      =   1'b0;
assign   tb_i_reset[263]                      =   1'b0;
assign   tb_i_sop[263]                        =   1'b0;
assign   tb_i_key_update[263]                 =   1'b0;
assign   tb_i_key[263]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[263]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[263]               =   1'b0;
assign   tb_i_rf_static_encrypt[263]          =   1'b1;
assign   tb_i_clear_fault_flags[263]          =   1'b0;
assign   tb_i_rf_static_aad_length[263]       =   64'h0000000000000100;
assign   tb_i_aad[263]                        =   tb_i_aad[262];
assign   tb_i_rf_static_plaintext_length[263] =   64'h0000000000000280;
assign   tb_i_plaintext[263]                  =   tb_i_plaintext[262];
assign   tb_o_valid[263]                      =   1'b0;
assign   tb_o_sop[263]                        =   1'b0;
assign   tb_o_ciphertext[263]                 =   tb_o_ciphertext[262];
assign   tb_o_tag_ready[263]                  =   1'b0;
assign   tb_o_tag[263]                        =   tb_o_tag[262];

// CLK no. 264/1240
// *************************************************
assign   tb_i_valid[264]                      =   1'b0;
assign   tb_i_reset[264]                      =   1'b0;
assign   tb_i_sop[264]                        =   1'b0;
assign   tb_i_key_update[264]                 =   1'b0;
assign   tb_i_key[264]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[264]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[264]               =   1'b0;
assign   tb_i_rf_static_encrypt[264]          =   1'b1;
assign   tb_i_clear_fault_flags[264]          =   1'b0;
assign   tb_i_rf_static_aad_length[264]       =   64'h0000000000000100;
assign   tb_i_aad[264]                        =   tb_i_aad[263];
assign   tb_i_rf_static_plaintext_length[264] =   64'h0000000000000280;
assign   tb_i_plaintext[264]                  =   tb_i_plaintext[263];
assign   tb_o_valid[264]                      =   1'b0;
assign   tb_o_sop[264]                        =   1'b0;
assign   tb_o_ciphertext[264]                 =   tb_o_ciphertext[263];
assign   tb_o_tag_ready[264]                  =   1'b0;
assign   tb_o_tag[264]                        =   tb_o_tag[263];

// CLK no. 265/1240
// *************************************************
assign   tb_i_valid[265]                      =   1'b0;
assign   tb_i_reset[265]                      =   1'b0;
assign   tb_i_sop[265]                        =   1'b0;
assign   tb_i_key_update[265]                 =   1'b0;
assign   tb_i_key[265]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[265]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[265]               =   1'b0;
assign   tb_i_rf_static_encrypt[265]          =   1'b1;
assign   tb_i_clear_fault_flags[265]          =   1'b0;
assign   tb_i_rf_static_aad_length[265]       =   64'h0000000000000100;
assign   tb_i_aad[265]                        =   tb_i_aad[264];
assign   tb_i_rf_static_plaintext_length[265] =   64'h0000000000000280;
assign   tb_i_plaintext[265]                  =   tb_i_plaintext[264];
assign   tb_o_valid[265]                      =   1'b0;
assign   tb_o_sop[265]                        =   1'b0;
assign   tb_o_ciphertext[265]                 =   tb_o_ciphertext[264];
assign   tb_o_tag_ready[265]                  =   1'b0;
assign   tb_o_tag[265]                        =   tb_o_tag[264];

// CLK no. 266/1240
// *************************************************
assign   tb_i_valid[266]                      =   1'b0;
assign   tb_i_reset[266]                      =   1'b0;
assign   tb_i_sop[266]                        =   1'b0;
assign   tb_i_key_update[266]                 =   1'b0;
assign   tb_i_key[266]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[266]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[266]               =   1'b0;
assign   tb_i_rf_static_encrypt[266]          =   1'b1;
assign   tb_i_clear_fault_flags[266]          =   1'b0;
assign   tb_i_rf_static_aad_length[266]       =   64'h0000000000000100;
assign   tb_i_aad[266]                        =   tb_i_aad[265];
assign   tb_i_rf_static_plaintext_length[266] =   64'h0000000000000280;
assign   tb_i_plaintext[266]                  =   tb_i_plaintext[265];
assign   tb_o_valid[266]                      =   1'b0;
assign   tb_o_sop[266]                        =   1'b0;
assign   tb_o_ciphertext[266]                 =   tb_o_ciphertext[265];
assign   tb_o_tag_ready[266]                  =   1'b0;
assign   tb_o_tag[266]                        =   tb_o_tag[265];

// CLK no. 267/1240
// *************************************************
assign   tb_i_valid[267]                      =   1'b0;
assign   tb_i_reset[267]                      =   1'b0;
assign   tb_i_sop[267]                        =   1'b0;
assign   tb_i_key_update[267]                 =   1'b0;
assign   tb_i_key[267]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[267]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[267]               =   1'b0;
assign   tb_i_rf_static_encrypt[267]          =   1'b1;
assign   tb_i_clear_fault_flags[267]          =   1'b0;
assign   tb_i_rf_static_aad_length[267]       =   64'h0000000000000100;
assign   tb_i_aad[267]                        =   tb_i_aad[266];
assign   tb_i_rf_static_plaintext_length[267] =   64'h0000000000000280;
assign   tb_i_plaintext[267]                  =   tb_i_plaintext[266];
assign   tb_o_valid[267]                      =   1'b0;
assign   tb_o_sop[267]                        =   1'b0;
assign   tb_o_ciphertext[267]                 =   tb_o_ciphertext[266];
assign   tb_o_tag_ready[267]                  =   1'b0;
assign   tb_o_tag[267]                        =   tb_o_tag[266];

// CLK no. 268/1240
// *************************************************
assign   tb_i_valid[268]                      =   1'b0;
assign   tb_i_reset[268]                      =   1'b0;
assign   tb_i_sop[268]                        =   1'b0;
assign   tb_i_key_update[268]                 =   1'b0;
assign   tb_i_key[268]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[268]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[268]               =   1'b0;
assign   tb_i_rf_static_encrypt[268]          =   1'b1;
assign   tb_i_clear_fault_flags[268]          =   1'b0;
assign   tb_i_rf_static_aad_length[268]       =   64'h0000000000000100;
assign   tb_i_aad[268]                        =   tb_i_aad[267];
assign   tb_i_rf_static_plaintext_length[268] =   64'h0000000000000280;
assign   tb_i_plaintext[268]                  =   tb_i_plaintext[267];
assign   tb_o_valid[268]                      =   1'b0;
assign   tb_o_sop[268]                        =   1'b0;
assign   tb_o_ciphertext[268]                 =   tb_o_ciphertext[267];
assign   tb_o_tag_ready[268]                  =   1'b0;
assign   tb_o_tag[268]                        =   tb_o_tag[267];

// CLK no. 269/1240
// *************************************************
assign   tb_i_valid[269]                      =   1'b0;
assign   tb_i_reset[269]                      =   1'b0;
assign   tb_i_sop[269]                        =   1'b0;
assign   tb_i_key_update[269]                 =   1'b0;
assign   tb_i_key[269]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[269]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[269]               =   1'b0;
assign   tb_i_rf_static_encrypt[269]          =   1'b1;
assign   tb_i_clear_fault_flags[269]          =   1'b0;
assign   tb_i_rf_static_aad_length[269]       =   64'h0000000000000100;
assign   tb_i_aad[269]                        =   tb_i_aad[268];
assign   tb_i_rf_static_plaintext_length[269] =   64'h0000000000000280;
assign   tb_i_plaintext[269]                  =   tb_i_plaintext[268];
assign   tb_o_valid[269]                      =   1'b0;
assign   tb_o_sop[269]                        =   1'b0;
assign   tb_o_ciphertext[269]                 =   tb_o_ciphertext[268];
assign   tb_o_tag_ready[269]                  =   1'b0;
assign   tb_o_tag[269]                        =   tb_o_tag[268];

// CLK no. 270/1240
// *************************************************
assign   tb_i_valid[270]                      =   1'b0;
assign   tb_i_reset[270]                      =   1'b0;
assign   tb_i_sop[270]                        =   1'b0;
assign   tb_i_key_update[270]                 =   1'b0;
assign   tb_i_key[270]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[270]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[270]               =   1'b0;
assign   tb_i_rf_static_encrypt[270]          =   1'b1;
assign   tb_i_clear_fault_flags[270]          =   1'b0;
assign   tb_i_rf_static_aad_length[270]       =   64'h0000000000000100;
assign   tb_i_aad[270]                        =   tb_i_aad[269];
assign   tb_i_rf_static_plaintext_length[270] =   64'h0000000000000280;
assign   tb_i_plaintext[270]                  =   tb_i_plaintext[269];
assign   tb_o_valid[270]                      =   1'b0;
assign   tb_o_sop[270]                        =   1'b0;
assign   tb_o_ciphertext[270]                 =   tb_o_ciphertext[269];
assign   tb_o_tag_ready[270]                  =   1'b0;
assign   tb_o_tag[270]                        =   tb_o_tag[269];

// CLK no. 271/1240
// *************************************************
assign   tb_i_valid[271]                      =   1'b0;
assign   tb_i_reset[271]                      =   1'b0;
assign   tb_i_sop[271]                        =   1'b0;
assign   tb_i_key_update[271]                 =   1'b0;
assign   tb_i_key[271]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[271]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[271]               =   1'b0;
assign   tb_i_rf_static_encrypt[271]          =   1'b1;
assign   tb_i_clear_fault_flags[271]          =   1'b0;
assign   tb_i_rf_static_aad_length[271]       =   64'h0000000000000100;
assign   tb_i_aad[271]                        =   tb_i_aad[270];
assign   tb_i_rf_static_plaintext_length[271] =   64'h0000000000000280;
assign   tb_i_plaintext[271]                  =   tb_i_plaintext[270];
assign   tb_o_valid[271]                      =   1'b0;
assign   tb_o_sop[271]                        =   1'b0;
assign   tb_o_ciphertext[271]                 =   tb_o_ciphertext[270];
assign   tb_o_tag_ready[271]                  =   1'b0;
assign   tb_o_tag[271]                        =   tb_o_tag[270];

// CLK no. 272/1240
// *************************************************
assign   tb_i_valid[272]                      =   1'b0;
assign   tb_i_reset[272]                      =   1'b0;
assign   tb_i_sop[272]                        =   1'b0;
assign   tb_i_key_update[272]                 =   1'b0;
assign   tb_i_key[272]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[272]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[272]               =   1'b0;
assign   tb_i_rf_static_encrypt[272]          =   1'b1;
assign   tb_i_clear_fault_flags[272]          =   1'b0;
assign   tb_i_rf_static_aad_length[272]       =   64'h0000000000000100;
assign   tb_i_aad[272]                        =   tb_i_aad[271];
assign   tb_i_rf_static_plaintext_length[272] =   64'h0000000000000280;
assign   tb_i_plaintext[272]                  =   tb_i_plaintext[271];
assign   tb_o_valid[272]                      =   1'b0;
assign   tb_o_sop[272]                        =   1'b0;
assign   tb_o_ciphertext[272]                 =   tb_o_ciphertext[271];
assign   tb_o_tag_ready[272]                  =   1'b0;
assign   tb_o_tag[272]                        =   tb_o_tag[271];

// CLK no. 273/1240
// *************************************************
assign   tb_i_valid[273]                      =   1'b0;
assign   tb_i_reset[273]                      =   1'b0;
assign   tb_i_sop[273]                        =   1'b0;
assign   tb_i_key_update[273]                 =   1'b0;
assign   tb_i_key[273]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[273]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[273]               =   1'b0;
assign   tb_i_rf_static_encrypt[273]          =   1'b1;
assign   tb_i_clear_fault_flags[273]          =   1'b0;
assign   tb_i_rf_static_aad_length[273]       =   64'h0000000000000100;
assign   tb_i_aad[273]                        =   tb_i_aad[272];
assign   tb_i_rf_static_plaintext_length[273] =   64'h0000000000000280;
assign   tb_i_plaintext[273]                  =   tb_i_plaintext[272];
assign   tb_o_valid[273]                      =   1'b0;
assign   tb_o_sop[273]                        =   1'b0;
assign   tb_o_ciphertext[273]                 =   tb_o_ciphertext[272];
assign   tb_o_tag_ready[273]                  =   1'b0;
assign   tb_o_tag[273]                        =   tb_o_tag[272];

// CLK no. 274/1240
// *************************************************
assign   tb_i_valid[274]                      =   1'b0;
assign   tb_i_reset[274]                      =   1'b0;
assign   tb_i_sop[274]                        =   1'b0;
assign   tb_i_key_update[274]                 =   1'b0;
assign   tb_i_key[274]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[274]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[274]               =   1'b0;
assign   tb_i_rf_static_encrypt[274]          =   1'b1;
assign   tb_i_clear_fault_flags[274]          =   1'b0;
assign   tb_i_rf_static_aad_length[274]       =   64'h0000000000000100;
assign   tb_i_aad[274]                        =   tb_i_aad[273];
assign   tb_i_rf_static_plaintext_length[274] =   64'h0000000000000280;
assign   tb_i_plaintext[274]                  =   tb_i_plaintext[273];
assign   tb_o_valid[274]                      =   1'b0;
assign   tb_o_sop[274]                        =   1'b0;
assign   tb_o_ciphertext[274]                 =   tb_o_ciphertext[273];
assign   tb_o_tag_ready[274]                  =   1'b0;
assign   tb_o_tag[274]                        =   tb_o_tag[273];

// CLK no. 275/1240
// *************************************************
assign   tb_i_valid[275]                      =   1'b0;
assign   tb_i_reset[275]                      =   1'b0;
assign   tb_i_sop[275]                        =   1'b0;
assign   tb_i_key_update[275]                 =   1'b0;
assign   tb_i_key[275]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[275]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[275]               =   1'b0;
assign   tb_i_rf_static_encrypt[275]          =   1'b1;
assign   tb_i_clear_fault_flags[275]          =   1'b0;
assign   tb_i_rf_static_aad_length[275]       =   64'h0000000000000100;
assign   tb_i_aad[275]                        =   tb_i_aad[274];
assign   tb_i_rf_static_plaintext_length[275] =   64'h0000000000000280;
assign   tb_i_plaintext[275]                  =   tb_i_plaintext[274];
assign   tb_o_valid[275]                      =   1'b0;
assign   tb_o_sop[275]                        =   1'b0;
assign   tb_o_ciphertext[275]                 =   tb_o_ciphertext[274];
assign   tb_o_tag_ready[275]                  =   1'b0;
assign   tb_o_tag[275]                        =   tb_o_tag[274];

// CLK no. 276/1240
// *************************************************
assign   tb_i_valid[276]                      =   1'b0;
assign   tb_i_reset[276]                      =   1'b0;
assign   tb_i_sop[276]                        =   1'b0;
assign   tb_i_key_update[276]                 =   1'b0;
assign   tb_i_key[276]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[276]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[276]               =   1'b0;
assign   tb_i_rf_static_encrypt[276]          =   1'b1;
assign   tb_i_clear_fault_flags[276]          =   1'b0;
assign   tb_i_rf_static_aad_length[276]       =   64'h0000000000000100;
assign   tb_i_aad[276]                        =   tb_i_aad[275];
assign   tb_i_rf_static_plaintext_length[276] =   64'h0000000000000280;
assign   tb_i_plaintext[276]                  =   tb_i_plaintext[275];
assign   tb_o_valid[276]                      =   1'b0;
assign   tb_o_sop[276]                        =   1'b0;
assign   tb_o_ciphertext[276]                 =   tb_o_ciphertext[275];
assign   tb_o_tag_ready[276]                  =   1'b0;
assign   tb_o_tag[276]                        =   tb_o_tag[275];

// CLK no. 277/1240
// *************************************************
assign   tb_i_valid[277]                      =   1'b0;
assign   tb_i_reset[277]                      =   1'b0;
assign   tb_i_sop[277]                        =   1'b0;
assign   tb_i_key_update[277]                 =   1'b0;
assign   tb_i_key[277]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[277]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[277]               =   1'b0;
assign   tb_i_rf_static_encrypt[277]          =   1'b1;
assign   tb_i_clear_fault_flags[277]          =   1'b0;
assign   tb_i_rf_static_aad_length[277]       =   64'h0000000000000100;
assign   tb_i_aad[277]                        =   tb_i_aad[276];
assign   tb_i_rf_static_plaintext_length[277] =   64'h0000000000000280;
assign   tb_i_plaintext[277]                  =   tb_i_plaintext[276];
assign   tb_o_valid[277]                      =   1'b0;
assign   tb_o_sop[277]                        =   1'b0;
assign   tb_o_ciphertext[277]                 =   tb_o_ciphertext[276];
assign   tb_o_tag_ready[277]                  =   1'b0;
assign   tb_o_tag[277]                        =   tb_o_tag[276];

// CLK no. 278/1240
// *************************************************
assign   tb_i_valid[278]                      =   1'b0;
assign   tb_i_reset[278]                      =   1'b0;
assign   tb_i_sop[278]                        =   1'b0;
assign   tb_i_key_update[278]                 =   1'b0;
assign   tb_i_key[278]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[278]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[278]               =   1'b0;
assign   tb_i_rf_static_encrypt[278]          =   1'b1;
assign   tb_i_clear_fault_flags[278]          =   1'b0;
assign   tb_i_rf_static_aad_length[278]       =   64'h0000000000000100;
assign   tb_i_aad[278]                        =   tb_i_aad[277];
assign   tb_i_rf_static_plaintext_length[278] =   64'h0000000000000280;
assign   tb_i_plaintext[278]                  =   tb_i_plaintext[277];
assign   tb_o_valid[278]                      =   1'b0;
assign   tb_o_sop[278]                        =   1'b0;
assign   tb_o_ciphertext[278]                 =   tb_o_ciphertext[277];
assign   tb_o_tag_ready[278]                  =   1'b0;
assign   tb_o_tag[278]                        =   tb_o_tag[277];

// CLK no. 279/1240
// *************************************************
assign   tb_i_valid[279]                      =   1'b0;
assign   tb_i_reset[279]                      =   1'b0;
assign   tb_i_sop[279]                        =   1'b0;
assign   tb_i_key_update[279]                 =   1'b0;
assign   tb_i_key[279]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[279]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[279]               =   1'b0;
assign   tb_i_rf_static_encrypt[279]          =   1'b1;
assign   tb_i_clear_fault_flags[279]          =   1'b0;
assign   tb_i_rf_static_aad_length[279]       =   64'h0000000000000100;
assign   tb_i_aad[279]                        =   tb_i_aad[278];
assign   tb_i_rf_static_plaintext_length[279] =   64'h0000000000000280;
assign   tb_i_plaintext[279]                  =   tb_i_plaintext[278];
assign   tb_o_valid[279]                      =   1'b0;
assign   tb_o_sop[279]                        =   1'b0;
assign   tb_o_ciphertext[279]                 =   tb_o_ciphertext[278];
assign   tb_o_tag_ready[279]                  =   1'b0;
assign   tb_o_tag[279]                        =   tb_o_tag[278];

// CLK no. 280/1240
// *************************************************
assign   tb_i_valid[280]                      =   1'b0;
assign   tb_i_reset[280]                      =   1'b0;
assign   tb_i_sop[280]                        =   1'b0;
assign   tb_i_key_update[280]                 =   1'b0;
assign   tb_i_key[280]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[280]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[280]               =   1'b0;
assign   tb_i_rf_static_encrypt[280]          =   1'b1;
assign   tb_i_clear_fault_flags[280]          =   1'b0;
assign   tb_i_rf_static_aad_length[280]       =   64'h0000000000000100;
assign   tb_i_aad[280]                        =   tb_i_aad[279];
assign   tb_i_rf_static_plaintext_length[280] =   64'h0000000000000280;
assign   tb_i_plaintext[280]                  =   tb_i_plaintext[279];
assign   tb_o_valid[280]                      =   1'b0;
assign   tb_o_sop[280]                        =   1'b0;
assign   tb_o_ciphertext[280]                 =   tb_o_ciphertext[279];
assign   tb_o_tag_ready[280]                  =   1'b0;
assign   tb_o_tag[280]                        =   tb_o_tag[279];

// CLK no. 281/1240
// *************************************************
assign   tb_i_valid[281]                      =   1'b0;
assign   tb_i_reset[281]                      =   1'b0;
assign   tb_i_sop[281]                        =   1'b0;
assign   tb_i_key_update[281]                 =   1'b0;
assign   tb_i_key[281]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[281]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[281]               =   1'b0;
assign   tb_i_rf_static_encrypt[281]          =   1'b1;
assign   tb_i_clear_fault_flags[281]          =   1'b0;
assign   tb_i_rf_static_aad_length[281]       =   64'h0000000000000100;
assign   tb_i_aad[281]                        =   tb_i_aad[280];
assign   tb_i_rf_static_plaintext_length[281] =   64'h0000000000000280;
assign   tb_i_plaintext[281]                  =   tb_i_plaintext[280];
assign   tb_o_valid[281]                      =   1'b0;
assign   tb_o_sop[281]                        =   1'b0;
assign   tb_o_ciphertext[281]                 =   tb_o_ciphertext[280];
assign   tb_o_tag_ready[281]                  =   1'b0;
assign   tb_o_tag[281]                        =   tb_o_tag[280];

// CLK no. 282/1240
// *************************************************
assign   tb_i_valid[282]                      =   1'b0;
assign   tb_i_reset[282]                      =   1'b0;
assign   tb_i_sop[282]                        =   1'b0;
assign   tb_i_key_update[282]                 =   1'b0;
assign   tb_i_key[282]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[282]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[282]               =   1'b0;
assign   tb_i_rf_static_encrypt[282]          =   1'b1;
assign   tb_i_clear_fault_flags[282]          =   1'b0;
assign   tb_i_rf_static_aad_length[282]       =   64'h0000000000000100;
assign   tb_i_aad[282]                        =   tb_i_aad[281];
assign   tb_i_rf_static_plaintext_length[282] =   64'h0000000000000280;
assign   tb_i_plaintext[282]                  =   tb_i_plaintext[281];
assign   tb_o_valid[282]                      =   1'b0;
assign   tb_o_sop[282]                        =   1'b0;
assign   tb_o_ciphertext[282]                 =   tb_o_ciphertext[281];
assign   tb_o_tag_ready[282]                  =   1'b0;
assign   tb_o_tag[282]                        =   tb_o_tag[281];

// CLK no. 283/1240
// *************************************************
assign   tb_i_valid[283]                      =   1'b0;
assign   tb_i_reset[283]                      =   1'b0;
assign   tb_i_sop[283]                        =   1'b0;
assign   tb_i_key_update[283]                 =   1'b0;
assign   tb_i_key[283]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[283]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[283]               =   1'b0;
assign   tb_i_rf_static_encrypt[283]          =   1'b1;
assign   tb_i_clear_fault_flags[283]          =   1'b0;
assign   tb_i_rf_static_aad_length[283]       =   64'h0000000000000100;
assign   tb_i_aad[283]                        =   tb_i_aad[282];
assign   tb_i_rf_static_plaintext_length[283] =   64'h0000000000000280;
assign   tb_i_plaintext[283]                  =   tb_i_plaintext[282];
assign   tb_o_valid[283]                      =   1'b1;
assign   tb_o_sop[283]                        =   1'b1;
assign   tb_o_ciphertext[283]                 =   256'h87f9b618fe00e02b852246d971002219e15ae94eb8b313ed489baac2e93f86a1;
assign   tb_o_tag_ready[283]                  =   1'b0;
assign   tb_o_tag[283]                        =   tb_o_tag[282];

// CLK no. 284/1240
// *************************************************
assign   tb_i_valid[284]                      =   1'b0;
assign   tb_i_reset[284]                      =   1'b0;
assign   tb_i_sop[284]                        =   1'b0;
assign   tb_i_key_update[284]                 =   1'b0;
assign   tb_i_key[284]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[284]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[284]               =   1'b0;
assign   tb_i_rf_static_encrypt[284]          =   1'b1;
assign   tb_i_clear_fault_flags[284]          =   1'b0;
assign   tb_i_rf_static_aad_length[284]       =   64'h0000000000000100;
assign   tb_i_aad[284]                        =   tb_i_aad[283];
assign   tb_i_rf_static_plaintext_length[284] =   64'h0000000000000280;
assign   tb_i_plaintext[284]                  =   tb_i_plaintext[283];
assign   tb_o_valid[284]                      =   1'b1;
assign   tb_o_sop[284]                        =   1'b0;
assign   tb_o_ciphertext[284]                 =   256'hcc291afe5735e94a00d241dec3d13f3e15a0caa283fb9ed6ee05618c58dc59a2;
assign   tb_o_tag_ready[284]                  =   1'b0;
assign   tb_o_tag[284]                        =   tb_o_tag[283];

// CLK no. 285/1240
// *************************************************
assign   tb_i_valid[285]                      =   1'b0;
assign   tb_i_reset[285]                      =   1'b0;
assign   tb_i_sop[285]                        =   1'b0;
assign   tb_i_key_update[285]                 =   1'b0;
assign   tb_i_key[285]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[285]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[285]               =   1'b0;
assign   tb_i_rf_static_encrypt[285]          =   1'b1;
assign   tb_i_clear_fault_flags[285]          =   1'b0;
assign   tb_i_rf_static_aad_length[285]       =   64'h0000000000000100;
assign   tb_i_aad[285]                        =   tb_i_aad[284];
assign   tb_i_rf_static_plaintext_length[285] =   64'h0000000000000280;
assign   tb_i_plaintext[285]                  =   tb_i_plaintext[284];
assign   tb_o_valid[285]                      =   1'b1;
assign   tb_o_sop[285]                        =   1'b0;
assign   tb_o_ciphertext[285]                 =   256'hd87b636884963a11709e140964a743b5;
assign   tb_o_tag_ready[285]                  =   1'b0;
assign   tb_o_tag[285]                        =   tb_o_tag[284];

// CLK no. 286/1240
// *************************************************
assign   tb_i_valid[286]                      =   1'b0;
assign   tb_i_reset[286]                      =   1'b0;
assign   tb_i_sop[286]                        =   1'b0;
assign   tb_i_key_update[286]                 =   1'b0;
assign   tb_i_key[286]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[286]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[286]               =   1'b0;
assign   tb_i_rf_static_encrypt[286]          =   1'b1;
assign   tb_i_clear_fault_flags[286]          =   1'b0;
assign   tb_i_rf_static_aad_length[286]       =   64'h0000000000000100;
assign   tb_i_aad[286]                        =   tb_i_aad[285];
assign   tb_i_rf_static_plaintext_length[286] =   64'h0000000000000280;
assign   tb_i_plaintext[286]                  =   tb_i_plaintext[285];
assign   tb_o_valid[286]                      =   1'b0;
assign   tb_o_sop[286]                        =   1'b0;
assign   tb_o_ciphertext[286]                 =   tb_o_ciphertext[285];
assign   tb_o_tag_ready[286]                  =   1'b0;
assign   tb_o_tag[286]                        =   tb_o_tag[285];

// CLK no. 287/1240
// *************************************************
assign   tb_i_valid[287]                      =   1'b0;
assign   tb_i_reset[287]                      =   1'b0;
assign   tb_i_sop[287]                        =   1'b0;
assign   tb_i_key_update[287]                 =   1'b0;
assign   tb_i_key[287]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[287]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[287]               =   1'b0;
assign   tb_i_rf_static_encrypt[287]          =   1'b1;
assign   tb_i_clear_fault_flags[287]          =   1'b0;
assign   tb_i_rf_static_aad_length[287]       =   64'h0000000000000100;
assign   tb_i_aad[287]                        =   tb_i_aad[286];
assign   tb_i_rf_static_plaintext_length[287] =   64'h0000000000000280;
assign   tb_i_plaintext[287]                  =   tb_i_plaintext[286];
assign   tb_o_valid[287]                      =   1'b0;
assign   tb_o_sop[287]                        =   1'b0;
assign   tb_o_ciphertext[287]                 =   tb_o_ciphertext[286];
assign   tb_o_tag_ready[287]                  =   1'b0;
assign   tb_o_tag[287]                        =   tb_o_tag[286];

// CLK no. 288/1240
// *************************************************
assign   tb_i_valid[288]                      =   1'b0;
assign   tb_i_reset[288]                      =   1'b0;
assign   tb_i_sop[288]                        =   1'b0;
assign   tb_i_key_update[288]                 =   1'b0;
assign   tb_i_key[288]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[288]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[288]               =   1'b0;
assign   tb_i_rf_static_encrypt[288]          =   1'b1;
assign   tb_i_clear_fault_flags[288]          =   1'b0;
assign   tb_i_rf_static_aad_length[288]       =   64'h0000000000000100;
assign   tb_i_aad[288]                        =   tb_i_aad[287];
assign   tb_i_rf_static_plaintext_length[288] =   64'h0000000000000280;
assign   tb_i_plaintext[288]                  =   tb_i_plaintext[287];
assign   tb_o_valid[288]                      =   1'b0;
assign   tb_o_sop[288]                        =   1'b0;
assign   tb_o_ciphertext[288]                 =   tb_o_ciphertext[287];
assign   tb_o_tag_ready[288]                  =   1'b0;
assign   tb_o_tag[288]                        =   tb_o_tag[287];

// CLK no. 289/1240
// *************************************************
assign   tb_i_valid[289]                      =   1'b0;
assign   tb_i_reset[289]                      =   1'b0;
assign   tb_i_sop[289]                        =   1'b0;
assign   tb_i_key_update[289]                 =   1'b0;
assign   tb_i_key[289]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[289]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[289]               =   1'b0;
assign   tb_i_rf_static_encrypt[289]          =   1'b1;
assign   tb_i_clear_fault_flags[289]          =   1'b0;
assign   tb_i_rf_static_aad_length[289]       =   64'h0000000000000100;
assign   tb_i_aad[289]                        =   tb_i_aad[288];
assign   tb_i_rf_static_plaintext_length[289] =   64'h0000000000000280;
assign   tb_i_plaintext[289]                  =   tb_i_plaintext[288];
assign   tb_o_valid[289]                      =   1'b0;
assign   tb_o_sop[289]                        =   1'b0;
assign   tb_o_ciphertext[289]                 =   tb_o_ciphertext[288];
assign   tb_o_tag_ready[289]                  =   1'b0;
assign   tb_o_tag[289]                        =   tb_o_tag[288];

// CLK no. 290/1240
// *************************************************
assign   tb_i_valid[290]                      =   1'b0;
assign   tb_i_reset[290]                      =   1'b0;
assign   tb_i_sop[290]                        =   1'b0;
assign   tb_i_key_update[290]                 =   1'b0;
assign   tb_i_key[290]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[290]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[290]               =   1'b0;
assign   tb_i_rf_static_encrypt[290]          =   1'b1;
assign   tb_i_clear_fault_flags[290]          =   1'b0;
assign   tb_i_rf_static_aad_length[290]       =   64'h0000000000000100;
assign   tb_i_aad[290]                        =   tb_i_aad[289];
assign   tb_i_rf_static_plaintext_length[290] =   64'h0000000000000280;
assign   tb_i_plaintext[290]                  =   tb_i_plaintext[289];
assign   tb_o_valid[290]                      =   1'b0;
assign   tb_o_sop[290]                        =   1'b0;
assign   tb_o_ciphertext[290]                 =   tb_o_ciphertext[289];
assign   tb_o_tag_ready[290]                  =   1'b0;
assign   tb_o_tag[290]                        =   tb_o_tag[289];

// CLK no. 291/1240
// *************************************************
assign   tb_i_valid[291]                      =   1'b0;
assign   tb_i_reset[291]                      =   1'b0;
assign   tb_i_sop[291]                        =   1'b0;
assign   tb_i_key_update[291]                 =   1'b0;
assign   tb_i_key[291]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[291]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[291]               =   1'b0;
assign   tb_i_rf_static_encrypt[291]          =   1'b1;
assign   tb_i_clear_fault_flags[291]          =   1'b0;
assign   tb_i_rf_static_aad_length[291]       =   64'h0000000000000100;
assign   tb_i_aad[291]                        =   tb_i_aad[290];
assign   tb_i_rf_static_plaintext_length[291] =   64'h0000000000000280;
assign   tb_i_plaintext[291]                  =   tb_i_plaintext[290];
assign   tb_o_valid[291]                      =   1'b0;
assign   tb_o_sop[291]                        =   1'b0;
assign   tb_o_ciphertext[291]                 =   tb_o_ciphertext[290];
assign   tb_o_tag_ready[291]                  =   1'b0;
assign   tb_o_tag[291]                        =   tb_o_tag[290];

// CLK no. 292/1240
// *************************************************
assign   tb_i_valid[292]                      =   1'b0;
assign   tb_i_reset[292]                      =   1'b0;
assign   tb_i_sop[292]                        =   1'b0;
assign   tb_i_key_update[292]                 =   1'b0;
assign   tb_i_key[292]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[292]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[292]               =   1'b0;
assign   tb_i_rf_static_encrypt[292]          =   1'b1;
assign   tb_i_clear_fault_flags[292]          =   1'b0;
assign   tb_i_rf_static_aad_length[292]       =   64'h0000000000000100;
assign   tb_i_aad[292]                        =   tb_i_aad[291];
assign   tb_i_rf_static_plaintext_length[292] =   64'h0000000000000280;
assign   tb_i_plaintext[292]                  =   tb_i_plaintext[291];
assign   tb_o_valid[292]                      =   1'b0;
assign   tb_o_sop[292]                        =   1'b0;
assign   tb_o_ciphertext[292]                 =   tb_o_ciphertext[291];
assign   tb_o_tag_ready[292]                  =   1'b0;
assign   tb_o_tag[292]                        =   tb_o_tag[291];

// CLK no. 293/1240
// *************************************************
assign   tb_i_valid[293]                      =   1'b0;
assign   tb_i_reset[293]                      =   1'b0;
assign   tb_i_sop[293]                        =   1'b0;
assign   tb_i_key_update[293]                 =   1'b0;
assign   tb_i_key[293]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[293]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[293]               =   1'b0;
assign   tb_i_rf_static_encrypt[293]          =   1'b1;
assign   tb_i_clear_fault_flags[293]          =   1'b0;
assign   tb_i_rf_static_aad_length[293]       =   64'h0000000000000100;
assign   tb_i_aad[293]                        =   tb_i_aad[292];
assign   tb_i_rf_static_plaintext_length[293] =   64'h0000000000000280;
assign   tb_i_plaintext[293]                  =   tb_i_plaintext[292];
assign   tb_o_valid[293]                      =   1'b0;
assign   tb_o_sop[293]                        =   1'b0;
assign   tb_o_ciphertext[293]                 =   tb_o_ciphertext[292];
assign   tb_o_tag_ready[293]                  =   1'b1;
assign   tb_o_tag[293]                        =   128'h8d691247d7fddc06d7ac0e6fd52d67bb;

// CLK no. 294/1240
// *************************************************
assign   tb_i_valid[294]                      =   1'b0;
assign   tb_i_reset[294]                      =   1'b0;
assign   tb_i_sop[294]                        =   1'b0;
assign   tb_i_key_update[294]                 =   1'b0;
assign   tb_i_key[294]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[294]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[294]               =   1'b0;
assign   tb_i_rf_static_encrypt[294]          =   1'b1;
assign   tb_i_clear_fault_flags[294]          =   1'b0;
assign   tb_i_rf_static_aad_length[294]       =   64'h0000000000000100;
assign   tb_i_aad[294]                        =   tb_i_aad[293];
assign   tb_i_rf_static_plaintext_length[294] =   64'h0000000000000280;
assign   tb_i_plaintext[294]                  =   tb_i_plaintext[293];
assign   tb_o_valid[294]                      =   1'b0;
assign   tb_o_sop[294]                        =   1'b0;
assign   tb_o_ciphertext[294]                 =   tb_o_ciphertext[293];
assign   tb_o_tag_ready[294]                  =   1'b0;
assign   tb_o_tag[294]                        =   tb_o_tag[293];

// CLK no. 295/1240
// *************************************************
assign   tb_i_valid[295]                      =   1'b0;
assign   tb_i_reset[295]                      =   1'b0;
assign   tb_i_sop[295]                        =   1'b0;
assign   tb_i_key_update[295]                 =   1'b0;
assign   tb_i_key[295]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[295]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[295]               =   1'b0;
assign   tb_i_rf_static_encrypt[295]          =   1'b1;
assign   tb_i_clear_fault_flags[295]          =   1'b0;
assign   tb_i_rf_static_aad_length[295]       =   64'h0000000000000100;
assign   tb_i_aad[295]                        =   tb_i_aad[294];
assign   tb_i_rf_static_plaintext_length[295] =   64'h0000000000000280;
assign   tb_i_plaintext[295]                  =   tb_i_plaintext[294];
assign   tb_o_valid[295]                      =   1'b0;
assign   tb_o_sop[295]                        =   1'b0;
assign   tb_o_ciphertext[295]                 =   tb_o_ciphertext[294];
assign   tb_o_tag_ready[295]                  =   1'b0;
assign   tb_o_tag[295]                        =   tb_o_tag[294];

// CLK no. 296/1240
// *************************************************
assign   tb_i_valid[296]                      =   1'b0;
assign   tb_i_reset[296]                      =   1'b0;
assign   tb_i_sop[296]                        =   1'b1;
assign   tb_i_key_update[296]                 =   1'b0;
assign   tb_i_key[296]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[296]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[296]               =   1'b0;
assign   tb_i_rf_static_encrypt[296]          =   1'b1;
assign   tb_i_clear_fault_flags[296]          =   1'b0;
assign   tb_i_rf_static_aad_length[296]       =   64'h0000000000000100;
assign   tb_i_aad[296]                        =   tb_i_aad[295];
assign   tb_i_rf_static_plaintext_length[296] =   64'h0000000000000280;
assign   tb_i_plaintext[296]                  =   tb_i_plaintext[295];
assign   tb_o_valid[296]                      =   1'b0;
assign   tb_o_sop[296]                        =   1'b0;
assign   tb_o_ciphertext[296]                 =   tb_o_ciphertext[295];
assign   tb_o_tag_ready[296]                  =   1'b0;
assign   tb_o_tag[296]                        =   tb_o_tag[295];

// CLK no. 297/1240
// *************************************************
assign   tb_i_valid[297]                      =   1'b1;
assign   tb_i_reset[297]                      =   1'b0;
assign   tb_i_sop[297]                        =   1'b0;
assign   tb_i_key_update[297]                 =   1'b0;
assign   tb_i_key[297]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[297]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[297]               =   1'b0;
assign   tb_i_rf_static_encrypt[297]          =   1'b1;
assign   tb_i_clear_fault_flags[297]          =   1'b0;
assign   tb_i_rf_static_aad_length[297]       =   64'h0000000000000100;
assign   tb_i_aad[297]                        =   256'h8e4b2d848cf4aac9a68fda26bb3c0eca8efbc1e30d59d3896758cb6213aa316b;
assign   tb_i_rf_static_plaintext_length[297] =   64'h0000000000000280;
assign   tb_i_plaintext[297]                  =   tb_i_plaintext[296];
assign   tb_o_valid[297]                      =   1'b0;
assign   tb_o_sop[297]                        =   1'b0;
assign   tb_o_ciphertext[297]                 =   tb_o_ciphertext[296];
assign   tb_o_tag_ready[297]                  =   1'b0;
assign   tb_o_tag[297]                        =   tb_o_tag[296];

// CLK no. 298/1240
// *************************************************
assign   tb_i_valid[298]                      =   1'b1;
assign   tb_i_reset[298]                      =   1'b0;
assign   tb_i_sop[298]                        =   1'b0;
assign   tb_i_key_update[298]                 =   1'b0;
assign   tb_i_key[298]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[298]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[298]               =   1'b0;
assign   tb_i_rf_static_encrypt[298]          =   1'b1;
assign   tb_i_clear_fault_flags[298]          =   1'b0;
assign   tb_i_rf_static_aad_length[298]       =   64'h0000000000000100;
assign   tb_i_aad[298]                        =   tb_i_aad[297];
assign   tb_i_rf_static_plaintext_length[298] =   64'h0000000000000280;
assign   tb_i_plaintext[298]                  =   256'h268cd4b32b1cff63c920c5074519bbfdb540a865cfcb12cf1d60ebff37e85ed1;
assign   tb_o_valid[298]                      =   1'b0;
assign   tb_o_sop[298]                        =   1'b0;
assign   tb_o_ciphertext[298]                 =   tb_o_ciphertext[297];
assign   tb_o_tag_ready[298]                  =   1'b0;
assign   tb_o_tag[298]                        =   tb_o_tag[297];

// CLK no. 299/1240
// *************************************************
assign   tb_i_valid[299]                      =   1'b1;
assign   tb_i_reset[299]                      =   1'b0;
assign   tb_i_sop[299]                        =   1'b0;
assign   tb_i_key_update[299]                 =   1'b0;
assign   tb_i_key[299]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[299]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[299]               =   1'b0;
assign   tb_i_rf_static_encrypt[299]          =   1'b1;
assign   tb_i_clear_fault_flags[299]          =   1'b0;
assign   tb_i_rf_static_aad_length[299]       =   64'h0000000000000100;
assign   tb_i_aad[299]                        =   tb_i_aad[298];
assign   tb_i_rf_static_plaintext_length[299] =   64'h0000000000000280;
assign   tb_i_plaintext[299]                  =   256'h372e6e63c1b7d9a99f82914e410ed1ae7a085beee5ef993e74a3c833ef6dde1d;
assign   tb_o_valid[299]                      =   1'b0;
assign   tb_o_sop[299]                        =   1'b0;
assign   tb_o_ciphertext[299]                 =   tb_o_ciphertext[298];
assign   tb_o_tag_ready[299]                  =   1'b0;
assign   tb_o_tag[299]                        =   tb_o_tag[298];

// CLK no. 300/1240
// *************************************************
assign   tb_i_valid[300]                      =   1'b1;
assign   tb_i_reset[300]                      =   1'b0;
assign   tb_i_sop[300]                        =   1'b0;
assign   tb_i_key_update[300]                 =   1'b0;
assign   tb_i_key[300]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[300]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[300]               =   1'b0;
assign   tb_i_rf_static_encrypt[300]          =   1'b1;
assign   tb_i_clear_fault_flags[300]          =   1'b0;
assign   tb_i_rf_static_aad_length[300]       =   64'h0000000000000100;
assign   tb_i_aad[300]                        =   tb_i_aad[299];
assign   tb_i_rf_static_plaintext_length[300] =   64'h0000000000000280;
assign   tb_i_plaintext[300]                  =   256'hf89e5041c8223c491ad7fc960b792e9f;
assign   tb_o_valid[300]                      =   1'b0;
assign   tb_o_sop[300]                        =   1'b0;
assign   tb_o_ciphertext[300]                 =   tb_o_ciphertext[299];
assign   tb_o_tag_ready[300]                  =   1'b0;
assign   tb_o_tag[300]                        =   tb_o_tag[299];

// CLK no. 301/1240
// *************************************************
assign   tb_i_valid[301]                      =   1'b0;
assign   tb_i_reset[301]                      =   1'b0;
assign   tb_i_sop[301]                        =   1'b0;
assign   tb_i_key_update[301]                 =   1'b0;
assign   tb_i_key[301]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[301]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[301]               =   1'b0;
assign   tb_i_rf_static_encrypt[301]          =   1'b1;
assign   tb_i_clear_fault_flags[301]          =   1'b0;
assign   tb_i_rf_static_aad_length[301]       =   64'h0000000000000100;
assign   tb_i_aad[301]                        =   tb_i_aad[300];
assign   tb_i_rf_static_plaintext_length[301] =   64'h0000000000000280;
assign   tb_i_plaintext[301]                  =   tb_i_plaintext[300];
assign   tb_o_valid[301]                      =   1'b0;
assign   tb_o_sop[301]                        =   1'b0;
assign   tb_o_ciphertext[301]                 =   tb_o_ciphertext[300];
assign   tb_o_tag_ready[301]                  =   1'b0;
assign   tb_o_tag[301]                        =   tb_o_tag[300];

// CLK no. 302/1240
// *************************************************
assign   tb_i_valid[302]                      =   1'b0;
assign   tb_i_reset[302]                      =   1'b0;
assign   tb_i_sop[302]                        =   1'b0;
assign   tb_i_key_update[302]                 =   1'b0;
assign   tb_i_key[302]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[302]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[302]               =   1'b0;
assign   tb_i_rf_static_encrypt[302]          =   1'b1;
assign   tb_i_clear_fault_flags[302]          =   1'b0;
assign   tb_i_rf_static_aad_length[302]       =   64'h0000000000000100;
assign   tb_i_aad[302]                        =   tb_i_aad[301];
assign   tb_i_rf_static_plaintext_length[302] =   64'h0000000000000280;
assign   tb_i_plaintext[302]                  =   tb_i_plaintext[301];
assign   tb_o_valid[302]                      =   1'b0;
assign   tb_o_sop[302]                        =   1'b0;
assign   tb_o_ciphertext[302]                 =   tb_o_ciphertext[301];
assign   tb_o_tag_ready[302]                  =   1'b0;
assign   tb_o_tag[302]                        =   tb_o_tag[301];

// CLK no. 303/1240
// *************************************************
assign   tb_i_valid[303]                      =   1'b0;
assign   tb_i_reset[303]                      =   1'b0;
assign   tb_i_sop[303]                        =   1'b0;
assign   tb_i_key_update[303]                 =   1'b0;
assign   tb_i_key[303]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[303]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[303]               =   1'b0;
assign   tb_i_rf_static_encrypt[303]          =   1'b1;
assign   tb_i_clear_fault_flags[303]          =   1'b0;
assign   tb_i_rf_static_aad_length[303]       =   64'h0000000000000100;
assign   tb_i_aad[303]                        =   tb_i_aad[302];
assign   tb_i_rf_static_plaintext_length[303] =   64'h0000000000000280;
assign   tb_i_plaintext[303]                  =   tb_i_plaintext[302];
assign   tb_o_valid[303]                      =   1'b0;
assign   tb_o_sop[303]                        =   1'b0;
assign   tb_o_ciphertext[303]                 =   tb_o_ciphertext[302];
assign   tb_o_tag_ready[303]                  =   1'b0;
assign   tb_o_tag[303]                        =   tb_o_tag[302];

// CLK no. 304/1240
// *************************************************
assign   tb_i_valid[304]                      =   1'b0;
assign   tb_i_reset[304]                      =   1'b0;
assign   tb_i_sop[304]                        =   1'b0;
assign   tb_i_key_update[304]                 =   1'b0;
assign   tb_i_key[304]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[304]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[304]               =   1'b0;
assign   tb_i_rf_static_encrypt[304]          =   1'b1;
assign   tb_i_clear_fault_flags[304]          =   1'b0;
assign   tb_i_rf_static_aad_length[304]       =   64'h0000000000000100;
assign   tb_i_aad[304]                        =   tb_i_aad[303];
assign   tb_i_rf_static_plaintext_length[304] =   64'h0000000000000280;
assign   tb_i_plaintext[304]                  =   tb_i_plaintext[303];
assign   tb_o_valid[304]                      =   1'b0;
assign   tb_o_sop[304]                        =   1'b0;
assign   tb_o_ciphertext[304]                 =   tb_o_ciphertext[303];
assign   tb_o_tag_ready[304]                  =   1'b0;
assign   tb_o_tag[304]                        =   tb_o_tag[303];

// CLK no. 305/1240
// *************************************************
assign   tb_i_valid[305]                      =   1'b0;
assign   tb_i_reset[305]                      =   1'b0;
assign   tb_i_sop[305]                        =   1'b0;
assign   tb_i_key_update[305]                 =   1'b0;
assign   tb_i_key[305]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[305]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[305]               =   1'b0;
assign   tb_i_rf_static_encrypt[305]          =   1'b1;
assign   tb_i_clear_fault_flags[305]          =   1'b0;
assign   tb_i_rf_static_aad_length[305]       =   64'h0000000000000100;
assign   tb_i_aad[305]                        =   tb_i_aad[304];
assign   tb_i_rf_static_plaintext_length[305] =   64'h0000000000000280;
assign   tb_i_plaintext[305]                  =   tb_i_plaintext[304];
assign   tb_o_valid[305]                      =   1'b0;
assign   tb_o_sop[305]                        =   1'b0;
assign   tb_o_ciphertext[305]                 =   tb_o_ciphertext[304];
assign   tb_o_tag_ready[305]                  =   1'b0;
assign   tb_o_tag[305]                        =   tb_o_tag[304];

// CLK no. 306/1240
// *************************************************
assign   tb_i_valid[306]                      =   1'b0;
assign   tb_i_reset[306]                      =   1'b0;
assign   tb_i_sop[306]                        =   1'b0;
assign   tb_i_key_update[306]                 =   1'b0;
assign   tb_i_key[306]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[306]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[306]               =   1'b0;
assign   tb_i_rf_static_encrypt[306]          =   1'b1;
assign   tb_i_clear_fault_flags[306]          =   1'b0;
assign   tb_i_rf_static_aad_length[306]       =   64'h0000000000000100;
assign   tb_i_aad[306]                        =   tb_i_aad[305];
assign   tb_i_rf_static_plaintext_length[306] =   64'h0000000000000280;
assign   tb_i_plaintext[306]                  =   tb_i_plaintext[305];
assign   tb_o_valid[306]                      =   1'b0;
assign   tb_o_sop[306]                        =   1'b0;
assign   tb_o_ciphertext[306]                 =   tb_o_ciphertext[305];
assign   tb_o_tag_ready[306]                  =   1'b0;
assign   tb_o_tag[306]                        =   tb_o_tag[305];

// CLK no. 307/1240
// *************************************************
assign   tb_i_valid[307]                      =   1'b0;
assign   tb_i_reset[307]                      =   1'b0;
assign   tb_i_sop[307]                        =   1'b0;
assign   tb_i_key_update[307]                 =   1'b0;
assign   tb_i_key[307]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[307]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[307]               =   1'b0;
assign   tb_i_rf_static_encrypt[307]          =   1'b1;
assign   tb_i_clear_fault_flags[307]          =   1'b0;
assign   tb_i_rf_static_aad_length[307]       =   64'h0000000000000100;
assign   tb_i_aad[307]                        =   tb_i_aad[306];
assign   tb_i_rf_static_plaintext_length[307] =   64'h0000000000000280;
assign   tb_i_plaintext[307]                  =   tb_i_plaintext[306];
assign   tb_o_valid[307]                      =   1'b0;
assign   tb_o_sop[307]                        =   1'b0;
assign   tb_o_ciphertext[307]                 =   tb_o_ciphertext[306];
assign   tb_o_tag_ready[307]                  =   1'b0;
assign   tb_o_tag[307]                        =   tb_o_tag[306];

// CLK no. 308/1240
// *************************************************
assign   tb_i_valid[308]                      =   1'b0;
assign   tb_i_reset[308]                      =   1'b0;
assign   tb_i_sop[308]                        =   1'b0;
assign   tb_i_key_update[308]                 =   1'b0;
assign   tb_i_key[308]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[308]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[308]               =   1'b0;
assign   tb_i_rf_static_encrypt[308]          =   1'b1;
assign   tb_i_clear_fault_flags[308]          =   1'b0;
assign   tb_i_rf_static_aad_length[308]       =   64'h0000000000000100;
assign   tb_i_aad[308]                        =   tb_i_aad[307];
assign   tb_i_rf_static_plaintext_length[308] =   64'h0000000000000280;
assign   tb_i_plaintext[308]                  =   tb_i_plaintext[307];
assign   tb_o_valid[308]                      =   1'b0;
assign   tb_o_sop[308]                        =   1'b0;
assign   tb_o_ciphertext[308]                 =   tb_o_ciphertext[307];
assign   tb_o_tag_ready[308]                  =   1'b0;
assign   tb_o_tag[308]                        =   tb_o_tag[307];

// CLK no. 309/1240
// *************************************************
assign   tb_i_valid[309]                      =   1'b0;
assign   tb_i_reset[309]                      =   1'b0;
assign   tb_i_sop[309]                        =   1'b0;
assign   tb_i_key_update[309]                 =   1'b0;
assign   tb_i_key[309]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[309]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[309]               =   1'b0;
assign   tb_i_rf_static_encrypt[309]          =   1'b1;
assign   tb_i_clear_fault_flags[309]          =   1'b0;
assign   tb_i_rf_static_aad_length[309]       =   64'h0000000000000100;
assign   tb_i_aad[309]                        =   tb_i_aad[308];
assign   tb_i_rf_static_plaintext_length[309] =   64'h0000000000000280;
assign   tb_i_plaintext[309]                  =   tb_i_plaintext[308];
assign   tb_o_valid[309]                      =   1'b0;
assign   tb_o_sop[309]                        =   1'b0;
assign   tb_o_ciphertext[309]                 =   tb_o_ciphertext[308];
assign   tb_o_tag_ready[309]                  =   1'b0;
assign   tb_o_tag[309]                        =   tb_o_tag[308];

// CLK no. 310/1240
// *************************************************
assign   tb_i_valid[310]                      =   1'b0;
assign   tb_i_reset[310]                      =   1'b0;
assign   tb_i_sop[310]                        =   1'b0;
assign   tb_i_key_update[310]                 =   1'b0;
assign   tb_i_key[310]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[310]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[310]               =   1'b0;
assign   tb_i_rf_static_encrypt[310]          =   1'b1;
assign   tb_i_clear_fault_flags[310]          =   1'b0;
assign   tb_i_rf_static_aad_length[310]       =   64'h0000000000000100;
assign   tb_i_aad[310]                        =   tb_i_aad[309];
assign   tb_i_rf_static_plaintext_length[310] =   64'h0000000000000280;
assign   tb_i_plaintext[310]                  =   tb_i_plaintext[309];
assign   tb_o_valid[310]                      =   1'b0;
assign   tb_o_sop[310]                        =   1'b0;
assign   tb_o_ciphertext[310]                 =   tb_o_ciphertext[309];
assign   tb_o_tag_ready[310]                  =   1'b0;
assign   tb_o_tag[310]                        =   tb_o_tag[309];

// CLK no. 311/1240
// *************************************************
assign   tb_i_valid[311]                      =   1'b0;
assign   tb_i_reset[311]                      =   1'b0;
assign   tb_i_sop[311]                        =   1'b0;
assign   tb_i_key_update[311]                 =   1'b0;
assign   tb_i_key[311]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[311]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[311]               =   1'b0;
assign   tb_i_rf_static_encrypt[311]          =   1'b1;
assign   tb_i_clear_fault_flags[311]          =   1'b0;
assign   tb_i_rf_static_aad_length[311]       =   64'h0000000000000100;
assign   tb_i_aad[311]                        =   tb_i_aad[310];
assign   tb_i_rf_static_plaintext_length[311] =   64'h0000000000000280;
assign   tb_i_plaintext[311]                  =   tb_i_plaintext[310];
assign   tb_o_valid[311]                      =   1'b0;
assign   tb_o_sop[311]                        =   1'b0;
assign   tb_o_ciphertext[311]                 =   tb_o_ciphertext[310];
assign   tb_o_tag_ready[311]                  =   1'b0;
assign   tb_o_tag[311]                        =   tb_o_tag[310];

// CLK no. 312/1240
// *************************************************
assign   tb_i_valid[312]                      =   1'b0;
assign   tb_i_reset[312]                      =   1'b0;
assign   tb_i_sop[312]                        =   1'b0;
assign   tb_i_key_update[312]                 =   1'b0;
assign   tb_i_key[312]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[312]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[312]               =   1'b0;
assign   tb_i_rf_static_encrypt[312]          =   1'b1;
assign   tb_i_clear_fault_flags[312]          =   1'b0;
assign   tb_i_rf_static_aad_length[312]       =   64'h0000000000000100;
assign   tb_i_aad[312]                        =   tb_i_aad[311];
assign   tb_i_rf_static_plaintext_length[312] =   64'h0000000000000280;
assign   tb_i_plaintext[312]                  =   tb_i_plaintext[311];
assign   tb_o_valid[312]                      =   1'b0;
assign   tb_o_sop[312]                        =   1'b0;
assign   tb_o_ciphertext[312]                 =   tb_o_ciphertext[311];
assign   tb_o_tag_ready[312]                  =   1'b0;
assign   tb_o_tag[312]                        =   tb_o_tag[311];

// CLK no. 313/1240
// *************************************************
assign   tb_i_valid[313]                      =   1'b0;
assign   tb_i_reset[313]                      =   1'b0;
assign   tb_i_sop[313]                        =   1'b0;
assign   tb_i_key_update[313]                 =   1'b0;
assign   tb_i_key[313]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[313]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[313]               =   1'b0;
assign   tb_i_rf_static_encrypt[313]          =   1'b1;
assign   tb_i_clear_fault_flags[313]          =   1'b0;
assign   tb_i_rf_static_aad_length[313]       =   64'h0000000000000100;
assign   tb_i_aad[313]                        =   tb_i_aad[312];
assign   tb_i_rf_static_plaintext_length[313] =   64'h0000000000000280;
assign   tb_i_plaintext[313]                  =   tb_i_plaintext[312];
assign   tb_o_valid[313]                      =   1'b0;
assign   tb_o_sop[313]                        =   1'b0;
assign   tb_o_ciphertext[313]                 =   tb_o_ciphertext[312];
assign   tb_o_tag_ready[313]                  =   1'b0;
assign   tb_o_tag[313]                        =   tb_o_tag[312];

// CLK no. 314/1240
// *************************************************
assign   tb_i_valid[314]                      =   1'b0;
assign   tb_i_reset[314]                      =   1'b0;
assign   tb_i_sop[314]                        =   1'b0;
assign   tb_i_key_update[314]                 =   1'b0;
assign   tb_i_key[314]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[314]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[314]               =   1'b0;
assign   tb_i_rf_static_encrypt[314]          =   1'b1;
assign   tb_i_clear_fault_flags[314]          =   1'b0;
assign   tb_i_rf_static_aad_length[314]       =   64'h0000000000000100;
assign   tb_i_aad[314]                        =   tb_i_aad[313];
assign   tb_i_rf_static_plaintext_length[314] =   64'h0000000000000280;
assign   tb_i_plaintext[314]                  =   tb_i_plaintext[313];
assign   tb_o_valid[314]                      =   1'b0;
assign   tb_o_sop[314]                        =   1'b0;
assign   tb_o_ciphertext[314]                 =   tb_o_ciphertext[313];
assign   tb_o_tag_ready[314]                  =   1'b0;
assign   tb_o_tag[314]                        =   tb_o_tag[313];

// CLK no. 315/1240
// *************************************************
assign   tb_i_valid[315]                      =   1'b0;
assign   tb_i_reset[315]                      =   1'b0;
assign   tb_i_sop[315]                        =   1'b0;
assign   tb_i_key_update[315]                 =   1'b0;
assign   tb_i_key[315]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[315]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[315]               =   1'b0;
assign   tb_i_rf_static_encrypt[315]          =   1'b1;
assign   tb_i_clear_fault_flags[315]          =   1'b0;
assign   tb_i_rf_static_aad_length[315]       =   64'h0000000000000100;
assign   tb_i_aad[315]                        =   tb_i_aad[314];
assign   tb_i_rf_static_plaintext_length[315] =   64'h0000000000000280;
assign   tb_i_plaintext[315]                  =   tb_i_plaintext[314];
assign   tb_o_valid[315]                      =   1'b0;
assign   tb_o_sop[315]                        =   1'b0;
assign   tb_o_ciphertext[315]                 =   tb_o_ciphertext[314];
assign   tb_o_tag_ready[315]                  =   1'b0;
assign   tb_o_tag[315]                        =   tb_o_tag[314];

// CLK no. 316/1240
// *************************************************
assign   tb_i_valid[316]                      =   1'b0;
assign   tb_i_reset[316]                      =   1'b0;
assign   tb_i_sop[316]                        =   1'b0;
assign   tb_i_key_update[316]                 =   1'b0;
assign   tb_i_key[316]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[316]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[316]               =   1'b0;
assign   tb_i_rf_static_encrypt[316]          =   1'b1;
assign   tb_i_clear_fault_flags[316]          =   1'b0;
assign   tb_i_rf_static_aad_length[316]       =   64'h0000000000000100;
assign   tb_i_aad[316]                        =   tb_i_aad[315];
assign   tb_i_rf_static_plaintext_length[316] =   64'h0000000000000280;
assign   tb_i_plaintext[316]                  =   tb_i_plaintext[315];
assign   tb_o_valid[316]                      =   1'b0;
assign   tb_o_sop[316]                        =   1'b0;
assign   tb_o_ciphertext[316]                 =   tb_o_ciphertext[315];
assign   tb_o_tag_ready[316]                  =   1'b0;
assign   tb_o_tag[316]                        =   tb_o_tag[315];

// CLK no. 317/1240
// *************************************************
assign   tb_i_valid[317]                      =   1'b0;
assign   tb_i_reset[317]                      =   1'b0;
assign   tb_i_sop[317]                        =   1'b0;
assign   tb_i_key_update[317]                 =   1'b0;
assign   tb_i_key[317]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[317]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[317]               =   1'b0;
assign   tb_i_rf_static_encrypt[317]          =   1'b1;
assign   tb_i_clear_fault_flags[317]          =   1'b0;
assign   tb_i_rf_static_aad_length[317]       =   64'h0000000000000100;
assign   tb_i_aad[317]                        =   tb_i_aad[316];
assign   tb_i_rf_static_plaintext_length[317] =   64'h0000000000000280;
assign   tb_i_plaintext[317]                  =   tb_i_plaintext[316];
assign   tb_o_valid[317]                      =   1'b0;
assign   tb_o_sop[317]                        =   1'b0;
assign   tb_o_ciphertext[317]                 =   tb_o_ciphertext[316];
assign   tb_o_tag_ready[317]                  =   1'b0;
assign   tb_o_tag[317]                        =   tb_o_tag[316];

// CLK no. 318/1240
// *************************************************
assign   tb_i_valid[318]                      =   1'b0;
assign   tb_i_reset[318]                      =   1'b0;
assign   tb_i_sop[318]                        =   1'b0;
assign   tb_i_key_update[318]                 =   1'b0;
assign   tb_i_key[318]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[318]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[318]               =   1'b0;
assign   tb_i_rf_static_encrypt[318]          =   1'b1;
assign   tb_i_clear_fault_flags[318]          =   1'b0;
assign   tb_i_rf_static_aad_length[318]       =   64'h0000000000000100;
assign   tb_i_aad[318]                        =   tb_i_aad[317];
assign   tb_i_rf_static_plaintext_length[318] =   64'h0000000000000280;
assign   tb_i_plaintext[318]                  =   tb_i_plaintext[317];
assign   tb_o_valid[318]                      =   1'b0;
assign   tb_o_sop[318]                        =   1'b0;
assign   tb_o_ciphertext[318]                 =   tb_o_ciphertext[317];
assign   tb_o_tag_ready[318]                  =   1'b0;
assign   tb_o_tag[318]                        =   tb_o_tag[317];

// CLK no. 319/1240
// *************************************************
assign   tb_i_valid[319]                      =   1'b0;
assign   tb_i_reset[319]                      =   1'b0;
assign   tb_i_sop[319]                        =   1'b0;
assign   tb_i_key_update[319]                 =   1'b0;
assign   tb_i_key[319]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[319]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[319]               =   1'b0;
assign   tb_i_rf_static_encrypt[319]          =   1'b1;
assign   tb_i_clear_fault_flags[319]          =   1'b0;
assign   tb_i_rf_static_aad_length[319]       =   64'h0000000000000100;
assign   tb_i_aad[319]                        =   tb_i_aad[318];
assign   tb_i_rf_static_plaintext_length[319] =   64'h0000000000000280;
assign   tb_i_plaintext[319]                  =   tb_i_plaintext[318];
assign   tb_o_valid[319]                      =   1'b0;
assign   tb_o_sop[319]                        =   1'b0;
assign   tb_o_ciphertext[319]                 =   tb_o_ciphertext[318];
assign   tb_o_tag_ready[319]                  =   1'b0;
assign   tb_o_tag[319]                        =   tb_o_tag[318];

// CLK no. 320/1240
// *************************************************
assign   tb_i_valid[320]                      =   1'b0;
assign   tb_i_reset[320]                      =   1'b0;
assign   tb_i_sop[320]                        =   1'b0;
assign   tb_i_key_update[320]                 =   1'b0;
assign   tb_i_key[320]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[320]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[320]               =   1'b0;
assign   tb_i_rf_static_encrypt[320]          =   1'b1;
assign   tb_i_clear_fault_flags[320]          =   1'b0;
assign   tb_i_rf_static_aad_length[320]       =   64'h0000000000000100;
assign   tb_i_aad[320]                        =   tb_i_aad[319];
assign   tb_i_rf_static_plaintext_length[320] =   64'h0000000000000280;
assign   tb_i_plaintext[320]                  =   tb_i_plaintext[319];
assign   tb_o_valid[320]                      =   1'b0;
assign   tb_o_sop[320]                        =   1'b0;
assign   tb_o_ciphertext[320]                 =   tb_o_ciphertext[319];
assign   tb_o_tag_ready[320]                  =   1'b0;
assign   tb_o_tag[320]                        =   tb_o_tag[319];

// CLK no. 321/1240
// *************************************************
assign   tb_i_valid[321]                      =   1'b0;
assign   tb_i_reset[321]                      =   1'b0;
assign   tb_i_sop[321]                        =   1'b0;
assign   tb_i_key_update[321]                 =   1'b0;
assign   tb_i_key[321]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[321]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[321]               =   1'b0;
assign   tb_i_rf_static_encrypt[321]          =   1'b1;
assign   tb_i_clear_fault_flags[321]          =   1'b0;
assign   tb_i_rf_static_aad_length[321]       =   64'h0000000000000100;
assign   tb_i_aad[321]                        =   tb_i_aad[320];
assign   tb_i_rf_static_plaintext_length[321] =   64'h0000000000000280;
assign   tb_i_plaintext[321]                  =   tb_i_plaintext[320];
assign   tb_o_valid[321]                      =   1'b0;
assign   tb_o_sop[321]                        =   1'b0;
assign   tb_o_ciphertext[321]                 =   tb_o_ciphertext[320];
assign   tb_o_tag_ready[321]                  =   1'b0;
assign   tb_o_tag[321]                        =   tb_o_tag[320];

// CLK no. 322/1240
// *************************************************
assign   tb_i_valid[322]                      =   1'b0;
assign   tb_i_reset[322]                      =   1'b0;
assign   tb_i_sop[322]                        =   1'b0;
assign   tb_i_key_update[322]                 =   1'b0;
assign   tb_i_key[322]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[322]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[322]               =   1'b0;
assign   tb_i_rf_static_encrypt[322]          =   1'b1;
assign   tb_i_clear_fault_flags[322]          =   1'b0;
assign   tb_i_rf_static_aad_length[322]       =   64'h0000000000000100;
assign   tb_i_aad[322]                        =   tb_i_aad[321];
assign   tb_i_rf_static_plaintext_length[322] =   64'h0000000000000280;
assign   tb_i_plaintext[322]                  =   tb_i_plaintext[321];
assign   tb_o_valid[322]                      =   1'b0;
assign   tb_o_sop[322]                        =   1'b0;
assign   tb_o_ciphertext[322]                 =   tb_o_ciphertext[321];
assign   tb_o_tag_ready[322]                  =   1'b0;
assign   tb_o_tag[322]                        =   tb_o_tag[321];

// CLK no. 323/1240
// *************************************************
assign   tb_i_valid[323]                      =   1'b0;
assign   tb_i_reset[323]                      =   1'b0;
assign   tb_i_sop[323]                        =   1'b0;
assign   tb_i_key_update[323]                 =   1'b0;
assign   tb_i_key[323]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[323]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[323]               =   1'b0;
assign   tb_i_rf_static_encrypt[323]          =   1'b1;
assign   tb_i_clear_fault_flags[323]          =   1'b0;
assign   tb_i_rf_static_aad_length[323]       =   64'h0000000000000100;
assign   tb_i_aad[323]                        =   tb_i_aad[322];
assign   tb_i_rf_static_plaintext_length[323] =   64'h0000000000000280;
assign   tb_i_plaintext[323]                  =   tb_i_plaintext[322];
assign   tb_o_valid[323]                      =   1'b0;
assign   tb_o_sop[323]                        =   1'b0;
assign   tb_o_ciphertext[323]                 =   tb_o_ciphertext[322];
assign   tb_o_tag_ready[323]                  =   1'b0;
assign   tb_o_tag[323]                        =   tb_o_tag[322];

// CLK no. 324/1240
// *************************************************
assign   tb_i_valid[324]                      =   1'b0;
assign   tb_i_reset[324]                      =   1'b0;
assign   tb_i_sop[324]                        =   1'b0;
assign   tb_i_key_update[324]                 =   1'b0;
assign   tb_i_key[324]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[324]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[324]               =   1'b0;
assign   tb_i_rf_static_encrypt[324]          =   1'b1;
assign   tb_i_clear_fault_flags[324]          =   1'b0;
assign   tb_i_rf_static_aad_length[324]       =   64'h0000000000000100;
assign   tb_i_aad[324]                        =   tb_i_aad[323];
assign   tb_i_rf_static_plaintext_length[324] =   64'h0000000000000280;
assign   tb_i_plaintext[324]                  =   tb_i_plaintext[323];
assign   tb_o_valid[324]                      =   1'b0;
assign   tb_o_sop[324]                        =   1'b0;
assign   tb_o_ciphertext[324]                 =   tb_o_ciphertext[323];
assign   tb_o_tag_ready[324]                  =   1'b0;
assign   tb_o_tag[324]                        =   tb_o_tag[323];

// CLK no. 325/1240
// *************************************************
assign   tb_i_valid[325]                      =   1'b0;
assign   tb_i_reset[325]                      =   1'b0;
assign   tb_i_sop[325]                        =   1'b0;
assign   tb_i_key_update[325]                 =   1'b0;
assign   tb_i_key[325]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[325]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[325]               =   1'b0;
assign   tb_i_rf_static_encrypt[325]          =   1'b1;
assign   tb_i_clear_fault_flags[325]          =   1'b0;
assign   tb_i_rf_static_aad_length[325]       =   64'h0000000000000100;
assign   tb_i_aad[325]                        =   tb_i_aad[324];
assign   tb_i_rf_static_plaintext_length[325] =   64'h0000000000000280;
assign   tb_i_plaintext[325]                  =   tb_i_plaintext[324];
assign   tb_o_valid[325]                      =   1'b0;
assign   tb_o_sop[325]                        =   1'b0;
assign   tb_o_ciphertext[325]                 =   tb_o_ciphertext[324];
assign   tb_o_tag_ready[325]                  =   1'b0;
assign   tb_o_tag[325]                        =   tb_o_tag[324];

// CLK no. 326/1240
// *************************************************
assign   tb_i_valid[326]                      =   1'b0;
assign   tb_i_reset[326]                      =   1'b0;
assign   tb_i_sop[326]                        =   1'b0;
assign   tb_i_key_update[326]                 =   1'b0;
assign   tb_i_key[326]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[326]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[326]               =   1'b0;
assign   tb_i_rf_static_encrypt[326]          =   1'b1;
assign   tb_i_clear_fault_flags[326]          =   1'b0;
assign   tb_i_rf_static_aad_length[326]       =   64'h0000000000000100;
assign   tb_i_aad[326]                        =   tb_i_aad[325];
assign   tb_i_rf_static_plaintext_length[326] =   64'h0000000000000280;
assign   tb_i_plaintext[326]                  =   tb_i_plaintext[325];
assign   tb_o_valid[326]                      =   1'b0;
assign   tb_o_sop[326]                        =   1'b0;
assign   tb_o_ciphertext[326]                 =   tb_o_ciphertext[325];
assign   tb_o_tag_ready[326]                  =   1'b0;
assign   tb_o_tag[326]                        =   tb_o_tag[325];

// CLK no. 327/1240
// *************************************************
assign   tb_i_valid[327]                      =   1'b0;
assign   tb_i_reset[327]                      =   1'b0;
assign   tb_i_sop[327]                        =   1'b0;
assign   tb_i_key_update[327]                 =   1'b0;
assign   tb_i_key[327]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[327]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[327]               =   1'b0;
assign   tb_i_rf_static_encrypt[327]          =   1'b1;
assign   tb_i_clear_fault_flags[327]          =   1'b0;
assign   tb_i_rf_static_aad_length[327]       =   64'h0000000000000100;
assign   tb_i_aad[327]                        =   tb_i_aad[326];
assign   tb_i_rf_static_plaintext_length[327] =   64'h0000000000000280;
assign   tb_i_plaintext[327]                  =   tb_i_plaintext[326];
assign   tb_o_valid[327]                      =   1'b0;
assign   tb_o_sop[327]                        =   1'b0;
assign   tb_o_ciphertext[327]                 =   tb_o_ciphertext[326];
assign   tb_o_tag_ready[327]                  =   1'b0;
assign   tb_o_tag[327]                        =   tb_o_tag[326];

// CLK no. 328/1240
// *************************************************
assign   tb_i_valid[328]                      =   1'b0;
assign   tb_i_reset[328]                      =   1'b0;
assign   tb_i_sop[328]                        =   1'b0;
assign   tb_i_key_update[328]                 =   1'b0;
assign   tb_i_key[328]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[328]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[328]               =   1'b0;
assign   tb_i_rf_static_encrypt[328]          =   1'b1;
assign   tb_i_clear_fault_flags[328]          =   1'b0;
assign   tb_i_rf_static_aad_length[328]       =   64'h0000000000000100;
assign   tb_i_aad[328]                        =   tb_i_aad[327];
assign   tb_i_rf_static_plaintext_length[328] =   64'h0000000000000280;
assign   tb_i_plaintext[328]                  =   tb_i_plaintext[327];
assign   tb_o_valid[328]                      =   1'b0;
assign   tb_o_sop[328]                        =   1'b0;
assign   tb_o_ciphertext[328]                 =   tb_o_ciphertext[327];
assign   tb_o_tag_ready[328]                  =   1'b0;
assign   tb_o_tag[328]                        =   tb_o_tag[327];

// CLK no. 329/1240
// *************************************************
assign   tb_i_valid[329]                      =   1'b0;
assign   tb_i_reset[329]                      =   1'b0;
assign   tb_i_sop[329]                        =   1'b0;
assign   tb_i_key_update[329]                 =   1'b0;
assign   tb_i_key[329]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[329]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[329]               =   1'b0;
assign   tb_i_rf_static_encrypt[329]          =   1'b1;
assign   tb_i_clear_fault_flags[329]          =   1'b0;
assign   tb_i_rf_static_aad_length[329]       =   64'h0000000000000100;
assign   tb_i_aad[329]                        =   tb_i_aad[328];
assign   tb_i_rf_static_plaintext_length[329] =   64'h0000000000000280;
assign   tb_i_plaintext[329]                  =   tb_i_plaintext[328];
assign   tb_o_valid[329]                      =   1'b0;
assign   tb_o_sop[329]                        =   1'b0;
assign   tb_o_ciphertext[329]                 =   tb_o_ciphertext[328];
assign   tb_o_tag_ready[329]                  =   1'b0;
assign   tb_o_tag[329]                        =   tb_o_tag[328];

// CLK no. 330/1240
// *************************************************
assign   tb_i_valid[330]                      =   1'b0;
assign   tb_i_reset[330]                      =   1'b0;
assign   tb_i_sop[330]                        =   1'b0;
assign   tb_i_key_update[330]                 =   1'b0;
assign   tb_i_key[330]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[330]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[330]               =   1'b0;
assign   tb_i_rf_static_encrypt[330]          =   1'b1;
assign   tb_i_clear_fault_flags[330]          =   1'b0;
assign   tb_i_rf_static_aad_length[330]       =   64'h0000000000000100;
assign   tb_i_aad[330]                        =   tb_i_aad[329];
assign   tb_i_rf_static_plaintext_length[330] =   64'h0000000000000280;
assign   tb_i_plaintext[330]                  =   tb_i_plaintext[329];
assign   tb_o_valid[330]                      =   1'b0;
assign   tb_o_sop[330]                        =   1'b0;
assign   tb_o_ciphertext[330]                 =   tb_o_ciphertext[329];
assign   tb_o_tag_ready[330]                  =   1'b0;
assign   tb_o_tag[330]                        =   tb_o_tag[329];

// CLK no. 331/1240
// *************************************************
assign   tb_i_valid[331]                      =   1'b0;
assign   tb_i_reset[331]                      =   1'b0;
assign   tb_i_sop[331]                        =   1'b0;
assign   tb_i_key_update[331]                 =   1'b0;
assign   tb_i_key[331]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[331]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[331]               =   1'b0;
assign   tb_i_rf_static_encrypt[331]          =   1'b1;
assign   tb_i_clear_fault_flags[331]          =   1'b0;
assign   tb_i_rf_static_aad_length[331]       =   64'h0000000000000100;
assign   tb_i_aad[331]                        =   tb_i_aad[330];
assign   tb_i_rf_static_plaintext_length[331] =   64'h0000000000000280;
assign   tb_i_plaintext[331]                  =   tb_i_plaintext[330];
assign   tb_o_valid[331]                      =   1'b0;
assign   tb_o_sop[331]                        =   1'b0;
assign   tb_o_ciphertext[331]                 =   tb_o_ciphertext[330];
assign   tb_o_tag_ready[331]                  =   1'b0;
assign   tb_o_tag[331]                        =   tb_o_tag[330];

// CLK no. 332/1240
// *************************************************
assign   tb_i_valid[332]                      =   1'b0;
assign   tb_i_reset[332]                      =   1'b0;
assign   tb_i_sop[332]                        =   1'b0;
assign   tb_i_key_update[332]                 =   1'b0;
assign   tb_i_key[332]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[332]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[332]               =   1'b0;
assign   tb_i_rf_static_encrypt[332]          =   1'b1;
assign   tb_i_clear_fault_flags[332]          =   1'b0;
assign   tb_i_rf_static_aad_length[332]       =   64'h0000000000000100;
assign   tb_i_aad[332]                        =   tb_i_aad[331];
assign   tb_i_rf_static_plaintext_length[332] =   64'h0000000000000280;
assign   tb_i_plaintext[332]                  =   tb_i_plaintext[331];
assign   tb_o_valid[332]                      =   1'b0;
assign   tb_o_sop[332]                        =   1'b0;
assign   tb_o_ciphertext[332]                 =   tb_o_ciphertext[331];
assign   tb_o_tag_ready[332]                  =   1'b0;
assign   tb_o_tag[332]                        =   tb_o_tag[331];

// CLK no. 333/1240
// *************************************************
assign   tb_i_valid[333]                      =   1'b0;
assign   tb_i_reset[333]                      =   1'b0;
assign   tb_i_sop[333]                        =   1'b0;
assign   tb_i_key_update[333]                 =   1'b0;
assign   tb_i_key[333]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[333]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[333]               =   1'b0;
assign   tb_i_rf_static_encrypt[333]          =   1'b1;
assign   tb_i_clear_fault_flags[333]          =   1'b0;
assign   tb_i_rf_static_aad_length[333]       =   64'h0000000000000100;
assign   tb_i_aad[333]                        =   tb_i_aad[332];
assign   tb_i_rf_static_plaintext_length[333] =   64'h0000000000000280;
assign   tb_i_plaintext[333]                  =   tb_i_plaintext[332];
assign   tb_o_valid[333]                      =   1'b0;
assign   tb_o_sop[333]                        =   1'b0;
assign   tb_o_ciphertext[333]                 =   tb_o_ciphertext[332];
assign   tb_o_tag_ready[333]                  =   1'b0;
assign   tb_o_tag[333]                        =   tb_o_tag[332];

// CLK no. 334/1240
// *************************************************
assign   tb_i_valid[334]                      =   1'b0;
assign   tb_i_reset[334]                      =   1'b0;
assign   tb_i_sop[334]                        =   1'b0;
assign   tb_i_key_update[334]                 =   1'b0;
assign   tb_i_key[334]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[334]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[334]               =   1'b0;
assign   tb_i_rf_static_encrypt[334]          =   1'b1;
assign   tb_i_clear_fault_flags[334]          =   1'b0;
assign   tb_i_rf_static_aad_length[334]       =   64'h0000000000000100;
assign   tb_i_aad[334]                        =   tb_i_aad[333];
assign   tb_i_rf_static_plaintext_length[334] =   64'h0000000000000280;
assign   tb_i_plaintext[334]                  =   tb_i_plaintext[333];
assign   tb_o_valid[334]                      =   1'b0;
assign   tb_o_sop[334]                        =   1'b0;
assign   tb_o_ciphertext[334]                 =   tb_o_ciphertext[333];
assign   tb_o_tag_ready[334]                  =   1'b0;
assign   tb_o_tag[334]                        =   tb_o_tag[333];

// CLK no. 335/1240
// *************************************************
assign   tb_i_valid[335]                      =   1'b0;
assign   tb_i_reset[335]                      =   1'b0;
assign   tb_i_sop[335]                        =   1'b0;
assign   tb_i_key_update[335]                 =   1'b0;
assign   tb_i_key[335]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[335]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[335]               =   1'b0;
assign   tb_i_rf_static_encrypt[335]          =   1'b1;
assign   tb_i_clear_fault_flags[335]          =   1'b0;
assign   tb_i_rf_static_aad_length[335]       =   64'h0000000000000100;
assign   tb_i_aad[335]                        =   tb_i_aad[334];
assign   tb_i_rf_static_plaintext_length[335] =   64'h0000000000000280;
assign   tb_i_plaintext[335]                  =   tb_i_plaintext[334];
assign   tb_o_valid[335]                      =   1'b0;
assign   tb_o_sop[335]                        =   1'b0;
assign   tb_o_ciphertext[335]                 =   tb_o_ciphertext[334];
assign   tb_o_tag_ready[335]                  =   1'b0;
assign   tb_o_tag[335]                        =   tb_o_tag[334];

// CLK no. 336/1240
// *************************************************
assign   tb_i_valid[336]                      =   1'b0;
assign   tb_i_reset[336]                      =   1'b0;
assign   tb_i_sop[336]                        =   1'b0;
assign   tb_i_key_update[336]                 =   1'b0;
assign   tb_i_key[336]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[336]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[336]               =   1'b0;
assign   tb_i_rf_static_encrypt[336]          =   1'b1;
assign   tb_i_clear_fault_flags[336]          =   1'b0;
assign   tb_i_rf_static_aad_length[336]       =   64'h0000000000000100;
assign   tb_i_aad[336]                        =   tb_i_aad[335];
assign   tb_i_rf_static_plaintext_length[336] =   64'h0000000000000280;
assign   tb_i_plaintext[336]                  =   tb_i_plaintext[335];
assign   tb_o_valid[336]                      =   1'b0;
assign   tb_o_sop[336]                        =   1'b0;
assign   tb_o_ciphertext[336]                 =   tb_o_ciphertext[335];
assign   tb_o_tag_ready[336]                  =   1'b0;
assign   tb_o_tag[336]                        =   tb_o_tag[335];

// CLK no. 337/1240
// *************************************************
assign   tb_i_valid[337]                      =   1'b0;
assign   tb_i_reset[337]                      =   1'b0;
assign   tb_i_sop[337]                        =   1'b0;
assign   tb_i_key_update[337]                 =   1'b0;
assign   tb_i_key[337]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[337]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[337]               =   1'b0;
assign   tb_i_rf_static_encrypt[337]          =   1'b1;
assign   tb_i_clear_fault_flags[337]          =   1'b0;
assign   tb_i_rf_static_aad_length[337]       =   64'h0000000000000100;
assign   tb_i_aad[337]                        =   tb_i_aad[336];
assign   tb_i_rf_static_plaintext_length[337] =   64'h0000000000000280;
assign   tb_i_plaintext[337]                  =   tb_i_plaintext[336];
assign   tb_o_valid[337]                      =   1'b0;
assign   tb_o_sop[337]                        =   1'b0;
assign   tb_o_ciphertext[337]                 =   tb_o_ciphertext[336];
assign   tb_o_tag_ready[337]                  =   1'b0;
assign   tb_o_tag[337]                        =   tb_o_tag[336];

// CLK no. 338/1240
// *************************************************
assign   tb_i_valid[338]                      =   1'b0;
assign   tb_i_reset[338]                      =   1'b0;
assign   tb_i_sop[338]                        =   1'b0;
assign   tb_i_key_update[338]                 =   1'b0;
assign   tb_i_key[338]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[338]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[338]               =   1'b0;
assign   tb_i_rf_static_encrypt[338]          =   1'b1;
assign   tb_i_clear_fault_flags[338]          =   1'b0;
assign   tb_i_rf_static_aad_length[338]       =   64'h0000000000000100;
assign   tb_i_aad[338]                        =   tb_i_aad[337];
assign   tb_i_rf_static_plaintext_length[338] =   64'h0000000000000280;
assign   tb_i_plaintext[338]                  =   tb_i_plaintext[337];
assign   tb_o_valid[338]                      =   1'b0;
assign   tb_o_sop[338]                        =   1'b0;
assign   tb_o_ciphertext[338]                 =   tb_o_ciphertext[337];
assign   tb_o_tag_ready[338]                  =   1'b0;
assign   tb_o_tag[338]                        =   tb_o_tag[337];

// CLK no. 339/1240
// *************************************************
assign   tb_i_valid[339]                      =   1'b0;
assign   tb_i_reset[339]                      =   1'b0;
assign   tb_i_sop[339]                        =   1'b0;
assign   tb_i_key_update[339]                 =   1'b0;
assign   tb_i_key[339]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[339]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[339]               =   1'b0;
assign   tb_i_rf_static_encrypt[339]          =   1'b1;
assign   tb_i_clear_fault_flags[339]          =   1'b0;
assign   tb_i_rf_static_aad_length[339]       =   64'h0000000000000100;
assign   tb_i_aad[339]                        =   tb_i_aad[338];
assign   tb_i_rf_static_plaintext_length[339] =   64'h0000000000000280;
assign   tb_i_plaintext[339]                  =   tb_i_plaintext[338];
assign   tb_o_valid[339]                      =   1'b0;
assign   tb_o_sop[339]                        =   1'b0;
assign   tb_o_ciphertext[339]                 =   tb_o_ciphertext[338];
assign   tb_o_tag_ready[339]                  =   1'b0;
assign   tb_o_tag[339]                        =   tb_o_tag[338];

// CLK no. 340/1240
// *************************************************
assign   tb_i_valid[340]                      =   1'b0;
assign   tb_i_reset[340]                      =   1'b0;
assign   tb_i_sop[340]                        =   1'b0;
assign   tb_i_key_update[340]                 =   1'b0;
assign   tb_i_key[340]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[340]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[340]               =   1'b0;
assign   tb_i_rf_static_encrypt[340]          =   1'b1;
assign   tb_i_clear_fault_flags[340]          =   1'b0;
assign   tb_i_rf_static_aad_length[340]       =   64'h0000000000000100;
assign   tb_i_aad[340]                        =   tb_i_aad[339];
assign   tb_i_rf_static_plaintext_length[340] =   64'h0000000000000280;
assign   tb_i_plaintext[340]                  =   tb_i_plaintext[339];
assign   tb_o_valid[340]                      =   1'b0;
assign   tb_o_sop[340]                        =   1'b0;
assign   tb_o_ciphertext[340]                 =   tb_o_ciphertext[339];
assign   tb_o_tag_ready[340]                  =   1'b0;
assign   tb_o_tag[340]                        =   tb_o_tag[339];

// CLK no. 341/1240
// *************************************************
assign   tb_i_valid[341]                      =   1'b0;
assign   tb_i_reset[341]                      =   1'b0;
assign   tb_i_sop[341]                        =   1'b0;
assign   tb_i_key_update[341]                 =   1'b0;
assign   tb_i_key[341]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[341]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[341]               =   1'b0;
assign   tb_i_rf_static_encrypt[341]          =   1'b1;
assign   tb_i_clear_fault_flags[341]          =   1'b0;
assign   tb_i_rf_static_aad_length[341]       =   64'h0000000000000100;
assign   tb_i_aad[341]                        =   tb_i_aad[340];
assign   tb_i_rf_static_plaintext_length[341] =   64'h0000000000000280;
assign   tb_i_plaintext[341]                  =   tb_i_plaintext[340];
assign   tb_o_valid[341]                      =   1'b0;
assign   tb_o_sop[341]                        =   1'b0;
assign   tb_o_ciphertext[341]                 =   tb_o_ciphertext[340];
assign   tb_o_tag_ready[341]                  =   1'b0;
assign   tb_o_tag[341]                        =   tb_o_tag[340];

// CLK no. 342/1240
// *************************************************
assign   tb_i_valid[342]                      =   1'b0;
assign   tb_i_reset[342]                      =   1'b0;
assign   tb_i_sop[342]                        =   1'b0;
assign   tb_i_key_update[342]                 =   1'b0;
assign   tb_i_key[342]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[342]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[342]               =   1'b0;
assign   tb_i_rf_static_encrypt[342]          =   1'b1;
assign   tb_i_clear_fault_flags[342]          =   1'b0;
assign   tb_i_rf_static_aad_length[342]       =   64'h0000000000000100;
assign   tb_i_aad[342]                        =   tb_i_aad[341];
assign   tb_i_rf_static_plaintext_length[342] =   64'h0000000000000280;
assign   tb_i_plaintext[342]                  =   tb_i_plaintext[341];
assign   tb_o_valid[342]                      =   1'b1;
assign   tb_o_sop[342]                        =   1'b1;
assign   tb_o_ciphertext[342]                 =   256'hc411f13c81cdc87092f45787ea7de0253e5c5bb0ae19692d4c46d599b2993a36;
assign   tb_o_tag_ready[342]                  =   1'b0;
assign   tb_o_tag[342]                        =   tb_o_tag[341];

// CLK no. 343/1240
// *************************************************
assign   tb_i_valid[343]                      =   1'b0;
assign   tb_i_reset[343]                      =   1'b0;
assign   tb_i_sop[343]                        =   1'b0;
assign   tb_i_key_update[343]                 =   1'b0;
assign   tb_i_key[343]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[343]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[343]               =   1'b0;
assign   tb_i_rf_static_encrypt[343]          =   1'b1;
assign   tb_i_clear_fault_flags[343]          =   1'b0;
assign   tb_i_rf_static_aad_length[343]       =   64'h0000000000000100;
assign   tb_i_aad[343]                        =   tb_i_aad[342];
assign   tb_i_rf_static_plaintext_length[343] =   64'h0000000000000280;
assign   tb_i_plaintext[343]                  =   tb_i_plaintext[342];
assign   tb_o_valid[343]                      =   1'b1;
assign   tb_o_sop[343]                        =   1'b0;
assign   tb_o_ciphertext[343]                 =   256'h43b29df5f80045f499281c15d2211656ea84d933298a2b50fcdc4d07f049e300;
assign   tb_o_tag_ready[343]                  =   1'b0;
assign   tb_o_tag[343]                        =   tb_o_tag[342];

// CLK no. 344/1240
// *************************************************
assign   tb_i_valid[344]                      =   1'b0;
assign   tb_i_reset[344]                      =   1'b0;
assign   tb_i_sop[344]                        =   1'b0;
assign   tb_i_key_update[344]                 =   1'b0;
assign   tb_i_key[344]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[344]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[344]               =   1'b0;
assign   tb_i_rf_static_encrypt[344]          =   1'b1;
assign   tb_i_clear_fault_flags[344]          =   1'b0;
assign   tb_i_rf_static_aad_length[344]       =   64'h0000000000000100;
assign   tb_i_aad[344]                        =   tb_i_aad[343];
assign   tb_i_rf_static_plaintext_length[344] =   64'h0000000000000280;
assign   tb_i_plaintext[344]                  =   tb_i_plaintext[343];
assign   tb_o_valid[344]                      =   1'b1;
assign   tb_o_sop[344]                        =   1'b0;
assign   tb_o_ciphertext[344]                 =   256'h9c312b1728cf41035242728bfd81ce70;
assign   tb_o_tag_ready[344]                  =   1'b0;
assign   tb_o_tag[344]                        =   tb_o_tag[343];

// CLK no. 345/1240
// *************************************************
assign   tb_i_valid[345]                      =   1'b0;
assign   tb_i_reset[345]                      =   1'b0;
assign   tb_i_sop[345]                        =   1'b0;
assign   tb_i_key_update[345]                 =   1'b0;
assign   tb_i_key[345]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[345]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[345]               =   1'b0;
assign   tb_i_rf_static_encrypt[345]          =   1'b1;
assign   tb_i_clear_fault_flags[345]          =   1'b0;
assign   tb_i_rf_static_aad_length[345]       =   64'h0000000000000100;
assign   tb_i_aad[345]                        =   tb_i_aad[344];
assign   tb_i_rf_static_plaintext_length[345] =   64'h0000000000000280;
assign   tb_i_plaintext[345]                  =   tb_i_plaintext[344];
assign   tb_o_valid[345]                      =   1'b0;
assign   tb_o_sop[345]                        =   1'b0;
assign   tb_o_ciphertext[345]                 =   tb_o_ciphertext[344];
assign   tb_o_tag_ready[345]                  =   1'b0;
assign   tb_o_tag[345]                        =   tb_o_tag[344];

// CLK no. 346/1240
// *************************************************
assign   tb_i_valid[346]                      =   1'b0;
assign   tb_i_reset[346]                      =   1'b0;
assign   tb_i_sop[346]                        =   1'b0;
assign   tb_i_key_update[346]                 =   1'b0;
assign   tb_i_key[346]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[346]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[346]               =   1'b0;
assign   tb_i_rf_static_encrypt[346]          =   1'b1;
assign   tb_i_clear_fault_flags[346]          =   1'b0;
assign   tb_i_rf_static_aad_length[346]       =   64'h0000000000000100;
assign   tb_i_aad[346]                        =   tb_i_aad[345];
assign   tb_i_rf_static_plaintext_length[346] =   64'h0000000000000280;
assign   tb_i_plaintext[346]                  =   tb_i_plaintext[345];
assign   tb_o_valid[346]                      =   1'b0;
assign   tb_o_sop[346]                        =   1'b0;
assign   tb_o_ciphertext[346]                 =   tb_o_ciphertext[345];
assign   tb_o_tag_ready[346]                  =   1'b0;
assign   tb_o_tag[346]                        =   tb_o_tag[345];

// CLK no. 347/1240
// *************************************************
assign   tb_i_valid[347]                      =   1'b0;
assign   tb_i_reset[347]                      =   1'b0;
assign   tb_i_sop[347]                        =   1'b0;
assign   tb_i_key_update[347]                 =   1'b0;
assign   tb_i_key[347]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[347]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[347]               =   1'b0;
assign   tb_i_rf_static_encrypt[347]          =   1'b1;
assign   tb_i_clear_fault_flags[347]          =   1'b0;
assign   tb_i_rf_static_aad_length[347]       =   64'h0000000000000100;
assign   tb_i_aad[347]                        =   tb_i_aad[346];
assign   tb_i_rf_static_plaintext_length[347] =   64'h0000000000000280;
assign   tb_i_plaintext[347]                  =   tb_i_plaintext[346];
assign   tb_o_valid[347]                      =   1'b0;
assign   tb_o_sop[347]                        =   1'b0;
assign   tb_o_ciphertext[347]                 =   tb_o_ciphertext[346];
assign   tb_o_tag_ready[347]                  =   1'b0;
assign   tb_o_tag[347]                        =   tb_o_tag[346];

// CLK no. 348/1240
// *************************************************
assign   tb_i_valid[348]                      =   1'b0;
assign   tb_i_reset[348]                      =   1'b0;
assign   tb_i_sop[348]                        =   1'b0;
assign   tb_i_key_update[348]                 =   1'b0;
assign   tb_i_key[348]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[348]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[348]               =   1'b0;
assign   tb_i_rf_static_encrypt[348]          =   1'b1;
assign   tb_i_clear_fault_flags[348]          =   1'b0;
assign   tb_i_rf_static_aad_length[348]       =   64'h0000000000000100;
assign   tb_i_aad[348]                        =   tb_i_aad[347];
assign   tb_i_rf_static_plaintext_length[348] =   64'h0000000000000280;
assign   tb_i_plaintext[348]                  =   tb_i_plaintext[347];
assign   tb_o_valid[348]                      =   1'b0;
assign   tb_o_sop[348]                        =   1'b0;
assign   tb_o_ciphertext[348]                 =   tb_o_ciphertext[347];
assign   tb_o_tag_ready[348]                  =   1'b0;
assign   tb_o_tag[348]                        =   tb_o_tag[347];

// CLK no. 349/1240
// *************************************************
assign   tb_i_valid[349]                      =   1'b0;
assign   tb_i_reset[349]                      =   1'b0;
assign   tb_i_sop[349]                        =   1'b0;
assign   tb_i_key_update[349]                 =   1'b0;
assign   tb_i_key[349]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[349]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[349]               =   1'b0;
assign   tb_i_rf_static_encrypt[349]          =   1'b1;
assign   tb_i_clear_fault_flags[349]          =   1'b0;
assign   tb_i_rf_static_aad_length[349]       =   64'h0000000000000100;
assign   tb_i_aad[349]                        =   tb_i_aad[348];
assign   tb_i_rf_static_plaintext_length[349] =   64'h0000000000000280;
assign   tb_i_plaintext[349]                  =   tb_i_plaintext[348];
assign   tb_o_valid[349]                      =   1'b0;
assign   tb_o_sop[349]                        =   1'b0;
assign   tb_o_ciphertext[349]                 =   tb_o_ciphertext[348];
assign   tb_o_tag_ready[349]                  =   1'b0;
assign   tb_o_tag[349]                        =   tb_o_tag[348];

// CLK no. 350/1240
// *************************************************
assign   tb_i_valid[350]                      =   1'b0;
assign   tb_i_reset[350]                      =   1'b0;
assign   tb_i_sop[350]                        =   1'b0;
assign   tb_i_key_update[350]                 =   1'b0;
assign   tb_i_key[350]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[350]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[350]               =   1'b0;
assign   tb_i_rf_static_encrypt[350]          =   1'b1;
assign   tb_i_clear_fault_flags[350]          =   1'b0;
assign   tb_i_rf_static_aad_length[350]       =   64'h0000000000000100;
assign   tb_i_aad[350]                        =   tb_i_aad[349];
assign   tb_i_rf_static_plaintext_length[350] =   64'h0000000000000280;
assign   tb_i_plaintext[350]                  =   tb_i_plaintext[349];
assign   tb_o_valid[350]                      =   1'b0;
assign   tb_o_sop[350]                        =   1'b0;
assign   tb_o_ciphertext[350]                 =   tb_o_ciphertext[349];
assign   tb_o_tag_ready[350]                  =   1'b0;
assign   tb_o_tag[350]                        =   tb_o_tag[349];

// CLK no. 351/1240
// *************************************************
assign   tb_i_valid[351]                      =   1'b0;
assign   tb_i_reset[351]                      =   1'b0;
assign   tb_i_sop[351]                        =   1'b0;
assign   tb_i_key_update[351]                 =   1'b0;
assign   tb_i_key[351]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[351]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[351]               =   1'b0;
assign   tb_i_rf_static_encrypt[351]          =   1'b1;
assign   tb_i_clear_fault_flags[351]          =   1'b0;
assign   tb_i_rf_static_aad_length[351]       =   64'h0000000000000100;
assign   tb_i_aad[351]                        =   tb_i_aad[350];
assign   tb_i_rf_static_plaintext_length[351] =   64'h0000000000000280;
assign   tb_i_plaintext[351]                  =   tb_i_plaintext[350];
assign   tb_o_valid[351]                      =   1'b0;
assign   tb_o_sop[351]                        =   1'b0;
assign   tb_o_ciphertext[351]                 =   tb_o_ciphertext[350];
assign   tb_o_tag_ready[351]                  =   1'b0;
assign   tb_o_tag[351]                        =   tb_o_tag[350];

// CLK no. 352/1240
// *************************************************
assign   tb_i_valid[352]                      =   1'b0;
assign   tb_i_reset[352]                      =   1'b0;
assign   tb_i_sop[352]                        =   1'b0;
assign   tb_i_key_update[352]                 =   1'b0;
assign   tb_i_key[352]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[352]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[352]               =   1'b0;
assign   tb_i_rf_static_encrypt[352]          =   1'b1;
assign   tb_i_clear_fault_flags[352]          =   1'b0;
assign   tb_i_rf_static_aad_length[352]       =   64'h0000000000000100;
assign   tb_i_aad[352]                        =   tb_i_aad[351];
assign   tb_i_rf_static_plaintext_length[352] =   64'h0000000000000280;
assign   tb_i_plaintext[352]                  =   tb_i_plaintext[351];
assign   tb_o_valid[352]                      =   1'b0;
assign   tb_o_sop[352]                        =   1'b0;
assign   tb_o_ciphertext[352]                 =   tb_o_ciphertext[351];
assign   tb_o_tag_ready[352]                  =   1'b1;
assign   tb_o_tag[352]                        =   128'h63aeab3b8d75b86848afb4c97ef9881f;

// CLK no. 353/1240
// *************************************************
assign   tb_i_valid[353]                      =   1'b0;
assign   tb_i_reset[353]                      =   1'b0;
assign   tb_i_sop[353]                        =   1'b0;
assign   tb_i_key_update[353]                 =   1'b0;
assign   tb_i_key[353]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[353]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[353]               =   1'b0;
assign   tb_i_rf_static_encrypt[353]          =   1'b1;
assign   tb_i_clear_fault_flags[353]          =   1'b0;
assign   tb_i_rf_static_aad_length[353]       =   64'h0000000000000100;
assign   tb_i_aad[353]                        =   tb_i_aad[352];
assign   tb_i_rf_static_plaintext_length[353] =   64'h0000000000000280;
assign   tb_i_plaintext[353]                  =   tb_i_plaintext[352];
assign   tb_o_valid[353]                      =   1'b0;
assign   tb_o_sop[353]                        =   1'b0;
assign   tb_o_ciphertext[353]                 =   tb_o_ciphertext[352];
assign   tb_o_tag_ready[353]                  =   1'b0;
assign   tb_o_tag[353]                        =   tb_o_tag[352];

// CLK no. 354/1240
// *************************************************
assign   tb_i_valid[354]                      =   1'b0;
assign   tb_i_reset[354]                      =   1'b0;
assign   tb_i_sop[354]                        =   1'b0;
assign   tb_i_key_update[354]                 =   1'b0;
assign   tb_i_key[354]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[354]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[354]               =   1'b0;
assign   tb_i_rf_static_encrypt[354]          =   1'b1;
assign   tb_i_clear_fault_flags[354]          =   1'b0;
assign   tb_i_rf_static_aad_length[354]       =   64'h0000000000000100;
assign   tb_i_aad[354]                        =   tb_i_aad[353];
assign   tb_i_rf_static_plaintext_length[354] =   64'h0000000000000280;
assign   tb_i_plaintext[354]                  =   tb_i_plaintext[353];
assign   tb_o_valid[354]                      =   1'b0;
assign   tb_o_sop[354]                        =   1'b0;
assign   tb_o_ciphertext[354]                 =   tb_o_ciphertext[353];
assign   tb_o_tag_ready[354]                  =   1'b0;
assign   tb_o_tag[354]                        =   tb_o_tag[353];

// CLK no. 355/1240
// *************************************************
assign   tb_i_valid[355]                      =   1'b0;
assign   tb_i_reset[355]                      =   1'b0;
assign   tb_i_sop[355]                        =   1'b1;
assign   tb_i_key_update[355]                 =   1'b0;
assign   tb_i_key[355]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[355]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[355]               =   1'b0;
assign   tb_i_rf_static_encrypt[355]          =   1'b1;
assign   tb_i_clear_fault_flags[355]          =   1'b0;
assign   tb_i_rf_static_aad_length[355]       =   64'h0000000000000100;
assign   tb_i_aad[355]                        =   tb_i_aad[354];
assign   tb_i_rf_static_plaintext_length[355] =   64'h0000000000000280;
assign   tb_i_plaintext[355]                  =   tb_i_plaintext[354];
assign   tb_o_valid[355]                      =   1'b0;
assign   tb_o_sop[355]                        =   1'b0;
assign   tb_o_ciphertext[355]                 =   tb_o_ciphertext[354];
assign   tb_o_tag_ready[355]                  =   1'b0;
assign   tb_o_tag[355]                        =   tb_o_tag[354];

// CLK no. 356/1240
// *************************************************
assign   tb_i_valid[356]                      =   1'b1;
assign   tb_i_reset[356]                      =   1'b0;
assign   tb_i_sop[356]                        =   1'b0;
assign   tb_i_key_update[356]                 =   1'b0;
assign   tb_i_key[356]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[356]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[356]               =   1'b0;
assign   tb_i_rf_static_encrypt[356]          =   1'b1;
assign   tb_i_clear_fault_flags[356]          =   1'b0;
assign   tb_i_rf_static_aad_length[356]       =   64'h0000000000000100;
assign   tb_i_aad[356]                        =   256'h6ba760801f42a697d8cacc28f47364609d20193e157a2b87b832141fb91df974;
assign   tb_i_rf_static_plaintext_length[356] =   64'h0000000000000280;
assign   tb_i_plaintext[356]                  =   tb_i_plaintext[355];
assign   tb_o_valid[356]                      =   1'b0;
assign   tb_o_sop[356]                        =   1'b0;
assign   tb_o_ciphertext[356]                 =   tb_o_ciphertext[355];
assign   tb_o_tag_ready[356]                  =   1'b0;
assign   tb_o_tag[356]                        =   tb_o_tag[355];

// CLK no. 357/1240
// *************************************************
assign   tb_i_valid[357]                      =   1'b1;
assign   tb_i_reset[357]                      =   1'b0;
assign   tb_i_sop[357]                        =   1'b0;
assign   tb_i_key_update[357]                 =   1'b0;
assign   tb_i_key[357]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[357]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[357]               =   1'b0;
assign   tb_i_rf_static_encrypt[357]          =   1'b1;
assign   tb_i_clear_fault_flags[357]          =   1'b0;
assign   tb_i_rf_static_aad_length[357]       =   64'h0000000000000100;
assign   tb_i_aad[357]                        =   tb_i_aad[356];
assign   tb_i_rf_static_plaintext_length[357] =   64'h0000000000000280;
assign   tb_i_plaintext[357]                  =   256'h1665676121ca4c012c59ffbb2f188236d572d59c01d250be47aeb4722a6b2166;
assign   tb_o_valid[357]                      =   1'b0;
assign   tb_o_sop[357]                        =   1'b0;
assign   tb_o_ciphertext[357]                 =   tb_o_ciphertext[356];
assign   tb_o_tag_ready[357]                  =   1'b0;
assign   tb_o_tag[357]                        =   tb_o_tag[356];

// CLK no. 358/1240
// *************************************************
assign   tb_i_valid[358]                      =   1'b1;
assign   tb_i_reset[358]                      =   1'b0;
assign   tb_i_sop[358]                        =   1'b0;
assign   tb_i_key_update[358]                 =   1'b0;
assign   tb_i_key[358]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[358]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[358]               =   1'b0;
assign   tb_i_rf_static_encrypt[358]          =   1'b1;
assign   tb_i_clear_fault_flags[358]          =   1'b0;
assign   tb_i_rf_static_aad_length[358]       =   64'h0000000000000100;
assign   tb_i_aad[358]                        =   tb_i_aad[357];
assign   tb_i_rf_static_plaintext_length[358] =   64'h0000000000000280;
assign   tb_i_plaintext[358]                  =   256'hadf959f7ecc5e9337342786cef3176ea40a44c607ed431a860a373201759cafd;
assign   tb_o_valid[358]                      =   1'b0;
assign   tb_o_sop[358]                        =   1'b0;
assign   tb_o_ciphertext[358]                 =   tb_o_ciphertext[357];
assign   tb_o_tag_ready[358]                  =   1'b0;
assign   tb_o_tag[358]                        =   tb_o_tag[357];

// CLK no. 359/1240
// *************************************************
assign   tb_i_valid[359]                      =   1'b1;
assign   tb_i_reset[359]                      =   1'b0;
assign   tb_i_sop[359]                        =   1'b0;
assign   tb_i_key_update[359]                 =   1'b0;
assign   tb_i_key[359]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[359]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[359]               =   1'b0;
assign   tb_i_rf_static_encrypt[359]          =   1'b1;
assign   tb_i_clear_fault_flags[359]          =   1'b0;
assign   tb_i_rf_static_aad_length[359]       =   64'h0000000000000100;
assign   tb_i_aad[359]                        =   tb_i_aad[358];
assign   tb_i_rf_static_plaintext_length[359] =   64'h0000000000000280;
assign   tb_i_plaintext[359]                  =   256'hc99de6c07b852df97be2061933961b7c;
assign   tb_o_valid[359]                      =   1'b0;
assign   tb_o_sop[359]                        =   1'b0;
assign   tb_o_ciphertext[359]                 =   tb_o_ciphertext[358];
assign   tb_o_tag_ready[359]                  =   1'b0;
assign   tb_o_tag[359]                        =   tb_o_tag[358];

// CLK no. 360/1240
// *************************************************
assign   tb_i_valid[360]                      =   1'b0;
assign   tb_i_reset[360]                      =   1'b0;
assign   tb_i_sop[360]                        =   1'b0;
assign   tb_i_key_update[360]                 =   1'b0;
assign   tb_i_key[360]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[360]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[360]               =   1'b0;
assign   tb_i_rf_static_encrypt[360]          =   1'b1;
assign   tb_i_clear_fault_flags[360]          =   1'b0;
assign   tb_i_rf_static_aad_length[360]       =   64'h0000000000000100;
assign   tb_i_aad[360]                        =   tb_i_aad[359];
assign   tb_i_rf_static_plaintext_length[360] =   64'h0000000000000280;
assign   tb_i_plaintext[360]                  =   tb_i_plaintext[359];
assign   tb_o_valid[360]                      =   1'b0;
assign   tb_o_sop[360]                        =   1'b0;
assign   tb_o_ciphertext[360]                 =   tb_o_ciphertext[359];
assign   tb_o_tag_ready[360]                  =   1'b0;
assign   tb_o_tag[360]                        =   tb_o_tag[359];

// CLK no. 361/1240
// *************************************************
assign   tb_i_valid[361]                      =   1'b0;
assign   tb_i_reset[361]                      =   1'b0;
assign   tb_i_sop[361]                        =   1'b0;
assign   tb_i_key_update[361]                 =   1'b0;
assign   tb_i_key[361]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[361]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[361]               =   1'b0;
assign   tb_i_rf_static_encrypt[361]          =   1'b1;
assign   tb_i_clear_fault_flags[361]          =   1'b0;
assign   tb_i_rf_static_aad_length[361]       =   64'h0000000000000100;
assign   tb_i_aad[361]                        =   tb_i_aad[360];
assign   tb_i_rf_static_plaintext_length[361] =   64'h0000000000000280;
assign   tb_i_plaintext[361]                  =   tb_i_plaintext[360];
assign   tb_o_valid[361]                      =   1'b0;
assign   tb_o_sop[361]                        =   1'b0;
assign   tb_o_ciphertext[361]                 =   tb_o_ciphertext[360];
assign   tb_o_tag_ready[361]                  =   1'b0;
assign   tb_o_tag[361]                        =   tb_o_tag[360];

// CLK no. 362/1240
// *************************************************
assign   tb_i_valid[362]                      =   1'b0;
assign   tb_i_reset[362]                      =   1'b0;
assign   tb_i_sop[362]                        =   1'b0;
assign   tb_i_key_update[362]                 =   1'b0;
assign   tb_i_key[362]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[362]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[362]               =   1'b0;
assign   tb_i_rf_static_encrypt[362]          =   1'b1;
assign   tb_i_clear_fault_flags[362]          =   1'b0;
assign   tb_i_rf_static_aad_length[362]       =   64'h0000000000000100;
assign   tb_i_aad[362]                        =   tb_i_aad[361];
assign   tb_i_rf_static_plaintext_length[362] =   64'h0000000000000280;
assign   tb_i_plaintext[362]                  =   tb_i_plaintext[361];
assign   tb_o_valid[362]                      =   1'b0;
assign   tb_o_sop[362]                        =   1'b0;
assign   tb_o_ciphertext[362]                 =   tb_o_ciphertext[361];
assign   tb_o_tag_ready[362]                  =   1'b0;
assign   tb_o_tag[362]                        =   tb_o_tag[361];

// CLK no. 363/1240
// *************************************************
assign   tb_i_valid[363]                      =   1'b0;
assign   tb_i_reset[363]                      =   1'b0;
assign   tb_i_sop[363]                        =   1'b0;
assign   tb_i_key_update[363]                 =   1'b0;
assign   tb_i_key[363]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[363]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[363]               =   1'b0;
assign   tb_i_rf_static_encrypt[363]          =   1'b1;
assign   tb_i_clear_fault_flags[363]          =   1'b0;
assign   tb_i_rf_static_aad_length[363]       =   64'h0000000000000100;
assign   tb_i_aad[363]                        =   tb_i_aad[362];
assign   tb_i_rf_static_plaintext_length[363] =   64'h0000000000000280;
assign   tb_i_plaintext[363]                  =   tb_i_plaintext[362];
assign   tb_o_valid[363]                      =   1'b0;
assign   tb_o_sop[363]                        =   1'b0;
assign   tb_o_ciphertext[363]                 =   tb_o_ciphertext[362];
assign   tb_o_tag_ready[363]                  =   1'b0;
assign   tb_o_tag[363]                        =   tb_o_tag[362];

// CLK no. 364/1240
// *************************************************
assign   tb_i_valid[364]                      =   1'b0;
assign   tb_i_reset[364]                      =   1'b0;
assign   tb_i_sop[364]                        =   1'b0;
assign   tb_i_key_update[364]                 =   1'b0;
assign   tb_i_key[364]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[364]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[364]               =   1'b0;
assign   tb_i_rf_static_encrypt[364]          =   1'b1;
assign   tb_i_clear_fault_flags[364]          =   1'b0;
assign   tb_i_rf_static_aad_length[364]       =   64'h0000000000000100;
assign   tb_i_aad[364]                        =   tb_i_aad[363];
assign   tb_i_rf_static_plaintext_length[364] =   64'h0000000000000280;
assign   tb_i_plaintext[364]                  =   tb_i_plaintext[363];
assign   tb_o_valid[364]                      =   1'b0;
assign   tb_o_sop[364]                        =   1'b0;
assign   tb_o_ciphertext[364]                 =   tb_o_ciphertext[363];
assign   tb_o_tag_ready[364]                  =   1'b0;
assign   tb_o_tag[364]                        =   tb_o_tag[363];

// CLK no. 365/1240
// *************************************************
assign   tb_i_valid[365]                      =   1'b0;
assign   tb_i_reset[365]                      =   1'b0;
assign   tb_i_sop[365]                        =   1'b0;
assign   tb_i_key_update[365]                 =   1'b0;
assign   tb_i_key[365]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[365]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[365]               =   1'b0;
assign   tb_i_rf_static_encrypt[365]          =   1'b1;
assign   tb_i_clear_fault_flags[365]          =   1'b0;
assign   tb_i_rf_static_aad_length[365]       =   64'h0000000000000100;
assign   tb_i_aad[365]                        =   tb_i_aad[364];
assign   tb_i_rf_static_plaintext_length[365] =   64'h0000000000000280;
assign   tb_i_plaintext[365]                  =   tb_i_plaintext[364];
assign   tb_o_valid[365]                      =   1'b0;
assign   tb_o_sop[365]                        =   1'b0;
assign   tb_o_ciphertext[365]                 =   tb_o_ciphertext[364];
assign   tb_o_tag_ready[365]                  =   1'b0;
assign   tb_o_tag[365]                        =   tb_o_tag[364];

// CLK no. 366/1240
// *************************************************
assign   tb_i_valid[366]                      =   1'b0;
assign   tb_i_reset[366]                      =   1'b0;
assign   tb_i_sop[366]                        =   1'b0;
assign   tb_i_key_update[366]                 =   1'b0;
assign   tb_i_key[366]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[366]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[366]               =   1'b0;
assign   tb_i_rf_static_encrypt[366]          =   1'b1;
assign   tb_i_clear_fault_flags[366]          =   1'b0;
assign   tb_i_rf_static_aad_length[366]       =   64'h0000000000000100;
assign   tb_i_aad[366]                        =   tb_i_aad[365];
assign   tb_i_rf_static_plaintext_length[366] =   64'h0000000000000280;
assign   tb_i_plaintext[366]                  =   tb_i_plaintext[365];
assign   tb_o_valid[366]                      =   1'b0;
assign   tb_o_sop[366]                        =   1'b0;
assign   tb_o_ciphertext[366]                 =   tb_o_ciphertext[365];
assign   tb_o_tag_ready[366]                  =   1'b0;
assign   tb_o_tag[366]                        =   tb_o_tag[365];

// CLK no. 367/1240
// *************************************************
assign   tb_i_valid[367]                      =   1'b0;
assign   tb_i_reset[367]                      =   1'b0;
assign   tb_i_sop[367]                        =   1'b0;
assign   tb_i_key_update[367]                 =   1'b0;
assign   tb_i_key[367]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[367]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[367]               =   1'b0;
assign   tb_i_rf_static_encrypt[367]          =   1'b1;
assign   tb_i_clear_fault_flags[367]          =   1'b0;
assign   tb_i_rf_static_aad_length[367]       =   64'h0000000000000100;
assign   tb_i_aad[367]                        =   tb_i_aad[366];
assign   tb_i_rf_static_plaintext_length[367] =   64'h0000000000000280;
assign   tb_i_plaintext[367]                  =   tb_i_plaintext[366];
assign   tb_o_valid[367]                      =   1'b0;
assign   tb_o_sop[367]                        =   1'b0;
assign   tb_o_ciphertext[367]                 =   tb_o_ciphertext[366];
assign   tb_o_tag_ready[367]                  =   1'b0;
assign   tb_o_tag[367]                        =   tb_o_tag[366];

// CLK no. 368/1240
// *************************************************
assign   tb_i_valid[368]                      =   1'b0;
assign   tb_i_reset[368]                      =   1'b0;
assign   tb_i_sop[368]                        =   1'b0;
assign   tb_i_key_update[368]                 =   1'b0;
assign   tb_i_key[368]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[368]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[368]               =   1'b0;
assign   tb_i_rf_static_encrypt[368]          =   1'b1;
assign   tb_i_clear_fault_flags[368]          =   1'b0;
assign   tb_i_rf_static_aad_length[368]       =   64'h0000000000000100;
assign   tb_i_aad[368]                        =   tb_i_aad[367];
assign   tb_i_rf_static_plaintext_length[368] =   64'h0000000000000280;
assign   tb_i_plaintext[368]                  =   tb_i_plaintext[367];
assign   tb_o_valid[368]                      =   1'b0;
assign   tb_o_sop[368]                        =   1'b0;
assign   tb_o_ciphertext[368]                 =   tb_o_ciphertext[367];
assign   tb_o_tag_ready[368]                  =   1'b0;
assign   tb_o_tag[368]                        =   tb_o_tag[367];

// CLK no. 369/1240
// *************************************************
assign   tb_i_valid[369]                      =   1'b0;
assign   tb_i_reset[369]                      =   1'b0;
assign   tb_i_sop[369]                        =   1'b0;
assign   tb_i_key_update[369]                 =   1'b0;
assign   tb_i_key[369]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[369]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[369]               =   1'b0;
assign   tb_i_rf_static_encrypt[369]          =   1'b1;
assign   tb_i_clear_fault_flags[369]          =   1'b0;
assign   tb_i_rf_static_aad_length[369]       =   64'h0000000000000100;
assign   tb_i_aad[369]                        =   tb_i_aad[368];
assign   tb_i_rf_static_plaintext_length[369] =   64'h0000000000000280;
assign   tb_i_plaintext[369]                  =   tb_i_plaintext[368];
assign   tb_o_valid[369]                      =   1'b0;
assign   tb_o_sop[369]                        =   1'b0;
assign   tb_o_ciphertext[369]                 =   tb_o_ciphertext[368];
assign   tb_o_tag_ready[369]                  =   1'b0;
assign   tb_o_tag[369]                        =   tb_o_tag[368];

// CLK no. 370/1240
// *************************************************
assign   tb_i_valid[370]                      =   1'b0;
assign   tb_i_reset[370]                      =   1'b0;
assign   tb_i_sop[370]                        =   1'b0;
assign   tb_i_key_update[370]                 =   1'b0;
assign   tb_i_key[370]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[370]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[370]               =   1'b0;
assign   tb_i_rf_static_encrypt[370]          =   1'b1;
assign   tb_i_clear_fault_flags[370]          =   1'b0;
assign   tb_i_rf_static_aad_length[370]       =   64'h0000000000000100;
assign   tb_i_aad[370]                        =   tb_i_aad[369];
assign   tb_i_rf_static_plaintext_length[370] =   64'h0000000000000280;
assign   tb_i_plaintext[370]                  =   tb_i_plaintext[369];
assign   tb_o_valid[370]                      =   1'b0;
assign   tb_o_sop[370]                        =   1'b0;
assign   tb_o_ciphertext[370]                 =   tb_o_ciphertext[369];
assign   tb_o_tag_ready[370]                  =   1'b0;
assign   tb_o_tag[370]                        =   tb_o_tag[369];

// CLK no. 371/1240
// *************************************************
assign   tb_i_valid[371]                      =   1'b0;
assign   tb_i_reset[371]                      =   1'b0;
assign   tb_i_sop[371]                        =   1'b0;
assign   tb_i_key_update[371]                 =   1'b0;
assign   tb_i_key[371]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[371]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[371]               =   1'b0;
assign   tb_i_rf_static_encrypt[371]          =   1'b1;
assign   tb_i_clear_fault_flags[371]          =   1'b0;
assign   tb_i_rf_static_aad_length[371]       =   64'h0000000000000100;
assign   tb_i_aad[371]                        =   tb_i_aad[370];
assign   tb_i_rf_static_plaintext_length[371] =   64'h0000000000000280;
assign   tb_i_plaintext[371]                  =   tb_i_plaintext[370];
assign   tb_o_valid[371]                      =   1'b0;
assign   tb_o_sop[371]                        =   1'b0;
assign   tb_o_ciphertext[371]                 =   tb_o_ciphertext[370];
assign   tb_o_tag_ready[371]                  =   1'b0;
assign   tb_o_tag[371]                        =   tb_o_tag[370];

// CLK no. 372/1240
// *************************************************
assign   tb_i_valid[372]                      =   1'b0;
assign   tb_i_reset[372]                      =   1'b0;
assign   tb_i_sop[372]                        =   1'b0;
assign   tb_i_key_update[372]                 =   1'b0;
assign   tb_i_key[372]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[372]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[372]               =   1'b0;
assign   tb_i_rf_static_encrypt[372]          =   1'b1;
assign   tb_i_clear_fault_flags[372]          =   1'b0;
assign   tb_i_rf_static_aad_length[372]       =   64'h0000000000000100;
assign   tb_i_aad[372]                        =   tb_i_aad[371];
assign   tb_i_rf_static_plaintext_length[372] =   64'h0000000000000280;
assign   tb_i_plaintext[372]                  =   tb_i_plaintext[371];
assign   tb_o_valid[372]                      =   1'b0;
assign   tb_o_sop[372]                        =   1'b0;
assign   tb_o_ciphertext[372]                 =   tb_o_ciphertext[371];
assign   tb_o_tag_ready[372]                  =   1'b0;
assign   tb_o_tag[372]                        =   tb_o_tag[371];

// CLK no. 373/1240
// *************************************************
assign   tb_i_valid[373]                      =   1'b0;
assign   tb_i_reset[373]                      =   1'b0;
assign   tb_i_sop[373]                        =   1'b0;
assign   tb_i_key_update[373]                 =   1'b0;
assign   tb_i_key[373]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[373]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[373]               =   1'b0;
assign   tb_i_rf_static_encrypt[373]          =   1'b1;
assign   tb_i_clear_fault_flags[373]          =   1'b0;
assign   tb_i_rf_static_aad_length[373]       =   64'h0000000000000100;
assign   tb_i_aad[373]                        =   tb_i_aad[372];
assign   tb_i_rf_static_plaintext_length[373] =   64'h0000000000000280;
assign   tb_i_plaintext[373]                  =   tb_i_plaintext[372];
assign   tb_o_valid[373]                      =   1'b0;
assign   tb_o_sop[373]                        =   1'b0;
assign   tb_o_ciphertext[373]                 =   tb_o_ciphertext[372];
assign   tb_o_tag_ready[373]                  =   1'b0;
assign   tb_o_tag[373]                        =   tb_o_tag[372];

// CLK no. 374/1240
// *************************************************
assign   tb_i_valid[374]                      =   1'b0;
assign   tb_i_reset[374]                      =   1'b0;
assign   tb_i_sop[374]                        =   1'b0;
assign   tb_i_key_update[374]                 =   1'b0;
assign   tb_i_key[374]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[374]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[374]               =   1'b0;
assign   tb_i_rf_static_encrypt[374]          =   1'b1;
assign   tb_i_clear_fault_flags[374]          =   1'b0;
assign   tb_i_rf_static_aad_length[374]       =   64'h0000000000000100;
assign   tb_i_aad[374]                        =   tb_i_aad[373];
assign   tb_i_rf_static_plaintext_length[374] =   64'h0000000000000280;
assign   tb_i_plaintext[374]                  =   tb_i_plaintext[373];
assign   tb_o_valid[374]                      =   1'b0;
assign   tb_o_sop[374]                        =   1'b0;
assign   tb_o_ciphertext[374]                 =   tb_o_ciphertext[373];
assign   tb_o_tag_ready[374]                  =   1'b0;
assign   tb_o_tag[374]                        =   tb_o_tag[373];

// CLK no. 375/1240
// *************************************************
assign   tb_i_valid[375]                      =   1'b0;
assign   tb_i_reset[375]                      =   1'b0;
assign   tb_i_sop[375]                        =   1'b0;
assign   tb_i_key_update[375]                 =   1'b0;
assign   tb_i_key[375]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[375]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[375]               =   1'b0;
assign   tb_i_rf_static_encrypt[375]          =   1'b1;
assign   tb_i_clear_fault_flags[375]          =   1'b0;
assign   tb_i_rf_static_aad_length[375]       =   64'h0000000000000100;
assign   tb_i_aad[375]                        =   tb_i_aad[374];
assign   tb_i_rf_static_plaintext_length[375] =   64'h0000000000000280;
assign   tb_i_plaintext[375]                  =   tb_i_plaintext[374];
assign   tb_o_valid[375]                      =   1'b0;
assign   tb_o_sop[375]                        =   1'b0;
assign   tb_o_ciphertext[375]                 =   tb_o_ciphertext[374];
assign   tb_o_tag_ready[375]                  =   1'b0;
assign   tb_o_tag[375]                        =   tb_o_tag[374];

// CLK no. 376/1240
// *************************************************
assign   tb_i_valid[376]                      =   1'b0;
assign   tb_i_reset[376]                      =   1'b0;
assign   tb_i_sop[376]                        =   1'b0;
assign   tb_i_key_update[376]                 =   1'b0;
assign   tb_i_key[376]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[376]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[376]               =   1'b0;
assign   tb_i_rf_static_encrypt[376]          =   1'b1;
assign   tb_i_clear_fault_flags[376]          =   1'b0;
assign   tb_i_rf_static_aad_length[376]       =   64'h0000000000000100;
assign   tb_i_aad[376]                        =   tb_i_aad[375];
assign   tb_i_rf_static_plaintext_length[376] =   64'h0000000000000280;
assign   tb_i_plaintext[376]                  =   tb_i_plaintext[375];
assign   tb_o_valid[376]                      =   1'b0;
assign   tb_o_sop[376]                        =   1'b0;
assign   tb_o_ciphertext[376]                 =   tb_o_ciphertext[375];
assign   tb_o_tag_ready[376]                  =   1'b0;
assign   tb_o_tag[376]                        =   tb_o_tag[375];

// CLK no. 377/1240
// *************************************************
assign   tb_i_valid[377]                      =   1'b0;
assign   tb_i_reset[377]                      =   1'b0;
assign   tb_i_sop[377]                        =   1'b0;
assign   tb_i_key_update[377]                 =   1'b0;
assign   tb_i_key[377]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[377]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[377]               =   1'b0;
assign   tb_i_rf_static_encrypt[377]          =   1'b1;
assign   tb_i_clear_fault_flags[377]          =   1'b0;
assign   tb_i_rf_static_aad_length[377]       =   64'h0000000000000100;
assign   tb_i_aad[377]                        =   tb_i_aad[376];
assign   tb_i_rf_static_plaintext_length[377] =   64'h0000000000000280;
assign   tb_i_plaintext[377]                  =   tb_i_plaintext[376];
assign   tb_o_valid[377]                      =   1'b0;
assign   tb_o_sop[377]                        =   1'b0;
assign   tb_o_ciphertext[377]                 =   tb_o_ciphertext[376];
assign   tb_o_tag_ready[377]                  =   1'b0;
assign   tb_o_tag[377]                        =   tb_o_tag[376];

// CLK no. 378/1240
// *************************************************
assign   tb_i_valid[378]                      =   1'b0;
assign   tb_i_reset[378]                      =   1'b0;
assign   tb_i_sop[378]                        =   1'b0;
assign   tb_i_key_update[378]                 =   1'b0;
assign   tb_i_key[378]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[378]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[378]               =   1'b0;
assign   tb_i_rf_static_encrypt[378]          =   1'b1;
assign   tb_i_clear_fault_flags[378]          =   1'b0;
assign   tb_i_rf_static_aad_length[378]       =   64'h0000000000000100;
assign   tb_i_aad[378]                        =   tb_i_aad[377];
assign   tb_i_rf_static_plaintext_length[378] =   64'h0000000000000280;
assign   tb_i_plaintext[378]                  =   tb_i_plaintext[377];
assign   tb_o_valid[378]                      =   1'b0;
assign   tb_o_sop[378]                        =   1'b0;
assign   tb_o_ciphertext[378]                 =   tb_o_ciphertext[377];
assign   tb_o_tag_ready[378]                  =   1'b0;
assign   tb_o_tag[378]                        =   tb_o_tag[377];

// CLK no. 379/1240
// *************************************************
assign   tb_i_valid[379]                      =   1'b0;
assign   tb_i_reset[379]                      =   1'b0;
assign   tb_i_sop[379]                        =   1'b0;
assign   tb_i_key_update[379]                 =   1'b0;
assign   tb_i_key[379]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[379]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[379]               =   1'b0;
assign   tb_i_rf_static_encrypt[379]          =   1'b1;
assign   tb_i_clear_fault_flags[379]          =   1'b0;
assign   tb_i_rf_static_aad_length[379]       =   64'h0000000000000100;
assign   tb_i_aad[379]                        =   tb_i_aad[378];
assign   tb_i_rf_static_plaintext_length[379] =   64'h0000000000000280;
assign   tb_i_plaintext[379]                  =   tb_i_plaintext[378];
assign   tb_o_valid[379]                      =   1'b0;
assign   tb_o_sop[379]                        =   1'b0;
assign   tb_o_ciphertext[379]                 =   tb_o_ciphertext[378];
assign   tb_o_tag_ready[379]                  =   1'b0;
assign   tb_o_tag[379]                        =   tb_o_tag[378];

// CLK no. 380/1240
// *************************************************
assign   tb_i_valid[380]                      =   1'b0;
assign   tb_i_reset[380]                      =   1'b0;
assign   tb_i_sop[380]                        =   1'b0;
assign   tb_i_key_update[380]                 =   1'b0;
assign   tb_i_key[380]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[380]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[380]               =   1'b0;
assign   tb_i_rf_static_encrypt[380]          =   1'b1;
assign   tb_i_clear_fault_flags[380]          =   1'b0;
assign   tb_i_rf_static_aad_length[380]       =   64'h0000000000000100;
assign   tb_i_aad[380]                        =   tb_i_aad[379];
assign   tb_i_rf_static_plaintext_length[380] =   64'h0000000000000280;
assign   tb_i_plaintext[380]                  =   tb_i_plaintext[379];
assign   tb_o_valid[380]                      =   1'b0;
assign   tb_o_sop[380]                        =   1'b0;
assign   tb_o_ciphertext[380]                 =   tb_o_ciphertext[379];
assign   tb_o_tag_ready[380]                  =   1'b0;
assign   tb_o_tag[380]                        =   tb_o_tag[379];

// CLK no. 381/1240
// *************************************************
assign   tb_i_valid[381]                      =   1'b0;
assign   tb_i_reset[381]                      =   1'b0;
assign   tb_i_sop[381]                        =   1'b0;
assign   tb_i_key_update[381]                 =   1'b0;
assign   tb_i_key[381]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[381]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[381]               =   1'b0;
assign   tb_i_rf_static_encrypt[381]          =   1'b1;
assign   tb_i_clear_fault_flags[381]          =   1'b0;
assign   tb_i_rf_static_aad_length[381]       =   64'h0000000000000100;
assign   tb_i_aad[381]                        =   tb_i_aad[380];
assign   tb_i_rf_static_plaintext_length[381] =   64'h0000000000000280;
assign   tb_i_plaintext[381]                  =   tb_i_plaintext[380];
assign   tb_o_valid[381]                      =   1'b0;
assign   tb_o_sop[381]                        =   1'b0;
assign   tb_o_ciphertext[381]                 =   tb_o_ciphertext[380];
assign   tb_o_tag_ready[381]                  =   1'b0;
assign   tb_o_tag[381]                        =   tb_o_tag[380];

// CLK no. 382/1240
// *************************************************
assign   tb_i_valid[382]                      =   1'b0;
assign   tb_i_reset[382]                      =   1'b0;
assign   tb_i_sop[382]                        =   1'b0;
assign   tb_i_key_update[382]                 =   1'b0;
assign   tb_i_key[382]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[382]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[382]               =   1'b0;
assign   tb_i_rf_static_encrypt[382]          =   1'b1;
assign   tb_i_clear_fault_flags[382]          =   1'b0;
assign   tb_i_rf_static_aad_length[382]       =   64'h0000000000000100;
assign   tb_i_aad[382]                        =   tb_i_aad[381];
assign   tb_i_rf_static_plaintext_length[382] =   64'h0000000000000280;
assign   tb_i_plaintext[382]                  =   tb_i_plaintext[381];
assign   tb_o_valid[382]                      =   1'b0;
assign   tb_o_sop[382]                        =   1'b0;
assign   tb_o_ciphertext[382]                 =   tb_o_ciphertext[381];
assign   tb_o_tag_ready[382]                  =   1'b0;
assign   tb_o_tag[382]                        =   tb_o_tag[381];

// CLK no. 383/1240
// *************************************************
assign   tb_i_valid[383]                      =   1'b0;
assign   tb_i_reset[383]                      =   1'b0;
assign   tb_i_sop[383]                        =   1'b0;
assign   tb_i_key_update[383]                 =   1'b0;
assign   tb_i_key[383]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[383]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[383]               =   1'b0;
assign   tb_i_rf_static_encrypt[383]          =   1'b1;
assign   tb_i_clear_fault_flags[383]          =   1'b0;
assign   tb_i_rf_static_aad_length[383]       =   64'h0000000000000100;
assign   tb_i_aad[383]                        =   tb_i_aad[382];
assign   tb_i_rf_static_plaintext_length[383] =   64'h0000000000000280;
assign   tb_i_plaintext[383]                  =   tb_i_plaintext[382];
assign   tb_o_valid[383]                      =   1'b0;
assign   tb_o_sop[383]                        =   1'b0;
assign   tb_o_ciphertext[383]                 =   tb_o_ciphertext[382];
assign   tb_o_tag_ready[383]                  =   1'b0;
assign   tb_o_tag[383]                        =   tb_o_tag[382];

// CLK no. 384/1240
// *************************************************
assign   tb_i_valid[384]                      =   1'b0;
assign   tb_i_reset[384]                      =   1'b0;
assign   tb_i_sop[384]                        =   1'b0;
assign   tb_i_key_update[384]                 =   1'b0;
assign   tb_i_key[384]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[384]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[384]               =   1'b0;
assign   tb_i_rf_static_encrypt[384]          =   1'b1;
assign   tb_i_clear_fault_flags[384]          =   1'b0;
assign   tb_i_rf_static_aad_length[384]       =   64'h0000000000000100;
assign   tb_i_aad[384]                        =   tb_i_aad[383];
assign   tb_i_rf_static_plaintext_length[384] =   64'h0000000000000280;
assign   tb_i_plaintext[384]                  =   tb_i_plaintext[383];
assign   tb_o_valid[384]                      =   1'b0;
assign   tb_o_sop[384]                        =   1'b0;
assign   tb_o_ciphertext[384]                 =   tb_o_ciphertext[383];
assign   tb_o_tag_ready[384]                  =   1'b0;
assign   tb_o_tag[384]                        =   tb_o_tag[383];

// CLK no. 385/1240
// *************************************************
assign   tb_i_valid[385]                      =   1'b0;
assign   tb_i_reset[385]                      =   1'b0;
assign   tb_i_sop[385]                        =   1'b0;
assign   tb_i_key_update[385]                 =   1'b0;
assign   tb_i_key[385]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[385]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[385]               =   1'b0;
assign   tb_i_rf_static_encrypt[385]          =   1'b1;
assign   tb_i_clear_fault_flags[385]          =   1'b0;
assign   tb_i_rf_static_aad_length[385]       =   64'h0000000000000100;
assign   tb_i_aad[385]                        =   tb_i_aad[384];
assign   tb_i_rf_static_plaintext_length[385] =   64'h0000000000000280;
assign   tb_i_plaintext[385]                  =   tb_i_plaintext[384];
assign   tb_o_valid[385]                      =   1'b0;
assign   tb_o_sop[385]                        =   1'b0;
assign   tb_o_ciphertext[385]                 =   tb_o_ciphertext[384];
assign   tb_o_tag_ready[385]                  =   1'b0;
assign   tb_o_tag[385]                        =   tb_o_tag[384];

// CLK no. 386/1240
// *************************************************
assign   tb_i_valid[386]                      =   1'b0;
assign   tb_i_reset[386]                      =   1'b0;
assign   tb_i_sop[386]                        =   1'b0;
assign   tb_i_key_update[386]                 =   1'b0;
assign   tb_i_key[386]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[386]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[386]               =   1'b0;
assign   tb_i_rf_static_encrypt[386]          =   1'b1;
assign   tb_i_clear_fault_flags[386]          =   1'b0;
assign   tb_i_rf_static_aad_length[386]       =   64'h0000000000000100;
assign   tb_i_aad[386]                        =   tb_i_aad[385];
assign   tb_i_rf_static_plaintext_length[386] =   64'h0000000000000280;
assign   tb_i_plaintext[386]                  =   tb_i_plaintext[385];
assign   tb_o_valid[386]                      =   1'b0;
assign   tb_o_sop[386]                        =   1'b0;
assign   tb_o_ciphertext[386]                 =   tb_o_ciphertext[385];
assign   tb_o_tag_ready[386]                  =   1'b0;
assign   tb_o_tag[386]                        =   tb_o_tag[385];

// CLK no. 387/1240
// *************************************************
assign   tb_i_valid[387]                      =   1'b0;
assign   tb_i_reset[387]                      =   1'b0;
assign   tb_i_sop[387]                        =   1'b0;
assign   tb_i_key_update[387]                 =   1'b0;
assign   tb_i_key[387]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[387]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[387]               =   1'b0;
assign   tb_i_rf_static_encrypt[387]          =   1'b1;
assign   tb_i_clear_fault_flags[387]          =   1'b0;
assign   tb_i_rf_static_aad_length[387]       =   64'h0000000000000100;
assign   tb_i_aad[387]                        =   tb_i_aad[386];
assign   tb_i_rf_static_plaintext_length[387] =   64'h0000000000000280;
assign   tb_i_plaintext[387]                  =   tb_i_plaintext[386];
assign   tb_o_valid[387]                      =   1'b0;
assign   tb_o_sop[387]                        =   1'b0;
assign   tb_o_ciphertext[387]                 =   tb_o_ciphertext[386];
assign   tb_o_tag_ready[387]                  =   1'b0;
assign   tb_o_tag[387]                        =   tb_o_tag[386];

// CLK no. 388/1240
// *************************************************
assign   tb_i_valid[388]                      =   1'b0;
assign   tb_i_reset[388]                      =   1'b0;
assign   tb_i_sop[388]                        =   1'b0;
assign   tb_i_key_update[388]                 =   1'b0;
assign   tb_i_key[388]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[388]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[388]               =   1'b0;
assign   tb_i_rf_static_encrypt[388]          =   1'b1;
assign   tb_i_clear_fault_flags[388]          =   1'b0;
assign   tb_i_rf_static_aad_length[388]       =   64'h0000000000000100;
assign   tb_i_aad[388]                        =   tb_i_aad[387];
assign   tb_i_rf_static_plaintext_length[388] =   64'h0000000000000280;
assign   tb_i_plaintext[388]                  =   tb_i_plaintext[387];
assign   tb_o_valid[388]                      =   1'b0;
assign   tb_o_sop[388]                        =   1'b0;
assign   tb_o_ciphertext[388]                 =   tb_o_ciphertext[387];
assign   tb_o_tag_ready[388]                  =   1'b0;
assign   tb_o_tag[388]                        =   tb_o_tag[387];

// CLK no. 389/1240
// *************************************************
assign   tb_i_valid[389]                      =   1'b0;
assign   tb_i_reset[389]                      =   1'b0;
assign   tb_i_sop[389]                        =   1'b0;
assign   tb_i_key_update[389]                 =   1'b0;
assign   tb_i_key[389]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[389]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[389]               =   1'b0;
assign   tb_i_rf_static_encrypt[389]          =   1'b1;
assign   tb_i_clear_fault_flags[389]          =   1'b0;
assign   tb_i_rf_static_aad_length[389]       =   64'h0000000000000100;
assign   tb_i_aad[389]                        =   tb_i_aad[388];
assign   tb_i_rf_static_plaintext_length[389] =   64'h0000000000000280;
assign   tb_i_plaintext[389]                  =   tb_i_plaintext[388];
assign   tb_o_valid[389]                      =   1'b0;
assign   tb_o_sop[389]                        =   1'b0;
assign   tb_o_ciphertext[389]                 =   tb_o_ciphertext[388];
assign   tb_o_tag_ready[389]                  =   1'b0;
assign   tb_o_tag[389]                        =   tb_o_tag[388];

// CLK no. 390/1240
// *************************************************
assign   tb_i_valid[390]                      =   1'b0;
assign   tb_i_reset[390]                      =   1'b0;
assign   tb_i_sop[390]                        =   1'b0;
assign   tb_i_key_update[390]                 =   1'b0;
assign   tb_i_key[390]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[390]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[390]               =   1'b0;
assign   tb_i_rf_static_encrypt[390]          =   1'b1;
assign   tb_i_clear_fault_flags[390]          =   1'b0;
assign   tb_i_rf_static_aad_length[390]       =   64'h0000000000000100;
assign   tb_i_aad[390]                        =   tb_i_aad[389];
assign   tb_i_rf_static_plaintext_length[390] =   64'h0000000000000280;
assign   tb_i_plaintext[390]                  =   tb_i_plaintext[389];
assign   tb_o_valid[390]                      =   1'b0;
assign   tb_o_sop[390]                        =   1'b0;
assign   tb_o_ciphertext[390]                 =   tb_o_ciphertext[389];
assign   tb_o_tag_ready[390]                  =   1'b0;
assign   tb_o_tag[390]                        =   tb_o_tag[389];

// CLK no. 391/1240
// *************************************************
assign   tb_i_valid[391]                      =   1'b0;
assign   tb_i_reset[391]                      =   1'b0;
assign   tb_i_sop[391]                        =   1'b0;
assign   tb_i_key_update[391]                 =   1'b0;
assign   tb_i_key[391]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[391]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[391]               =   1'b0;
assign   tb_i_rf_static_encrypt[391]          =   1'b1;
assign   tb_i_clear_fault_flags[391]          =   1'b0;
assign   tb_i_rf_static_aad_length[391]       =   64'h0000000000000100;
assign   tb_i_aad[391]                        =   tb_i_aad[390];
assign   tb_i_rf_static_plaintext_length[391] =   64'h0000000000000280;
assign   tb_i_plaintext[391]                  =   tb_i_plaintext[390];
assign   tb_o_valid[391]                      =   1'b0;
assign   tb_o_sop[391]                        =   1'b0;
assign   tb_o_ciphertext[391]                 =   tb_o_ciphertext[390];
assign   tb_o_tag_ready[391]                  =   1'b0;
assign   tb_o_tag[391]                        =   tb_o_tag[390];

// CLK no. 392/1240
// *************************************************
assign   tb_i_valid[392]                      =   1'b0;
assign   tb_i_reset[392]                      =   1'b0;
assign   tb_i_sop[392]                        =   1'b0;
assign   tb_i_key_update[392]                 =   1'b0;
assign   tb_i_key[392]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[392]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[392]               =   1'b0;
assign   tb_i_rf_static_encrypt[392]          =   1'b1;
assign   tb_i_clear_fault_flags[392]          =   1'b0;
assign   tb_i_rf_static_aad_length[392]       =   64'h0000000000000100;
assign   tb_i_aad[392]                        =   tb_i_aad[391];
assign   tb_i_rf_static_plaintext_length[392] =   64'h0000000000000280;
assign   tb_i_plaintext[392]                  =   tb_i_plaintext[391];
assign   tb_o_valid[392]                      =   1'b0;
assign   tb_o_sop[392]                        =   1'b0;
assign   tb_o_ciphertext[392]                 =   tb_o_ciphertext[391];
assign   tb_o_tag_ready[392]                  =   1'b0;
assign   tb_o_tag[392]                        =   tb_o_tag[391];

// CLK no. 393/1240
// *************************************************
assign   tb_i_valid[393]                      =   1'b0;
assign   tb_i_reset[393]                      =   1'b0;
assign   tb_i_sop[393]                        =   1'b0;
assign   tb_i_key_update[393]                 =   1'b0;
assign   tb_i_key[393]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[393]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[393]               =   1'b0;
assign   tb_i_rf_static_encrypt[393]          =   1'b1;
assign   tb_i_clear_fault_flags[393]          =   1'b0;
assign   tb_i_rf_static_aad_length[393]       =   64'h0000000000000100;
assign   tb_i_aad[393]                        =   tb_i_aad[392];
assign   tb_i_rf_static_plaintext_length[393] =   64'h0000000000000280;
assign   tb_i_plaintext[393]                  =   tb_i_plaintext[392];
assign   tb_o_valid[393]                      =   1'b0;
assign   tb_o_sop[393]                        =   1'b0;
assign   tb_o_ciphertext[393]                 =   tb_o_ciphertext[392];
assign   tb_o_tag_ready[393]                  =   1'b0;
assign   tb_o_tag[393]                        =   tb_o_tag[392];

// CLK no. 394/1240
// *************************************************
assign   tb_i_valid[394]                      =   1'b0;
assign   tb_i_reset[394]                      =   1'b0;
assign   tb_i_sop[394]                        =   1'b0;
assign   tb_i_key_update[394]                 =   1'b0;
assign   tb_i_key[394]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[394]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[394]               =   1'b0;
assign   tb_i_rf_static_encrypt[394]          =   1'b1;
assign   tb_i_clear_fault_flags[394]          =   1'b0;
assign   tb_i_rf_static_aad_length[394]       =   64'h0000000000000100;
assign   tb_i_aad[394]                        =   tb_i_aad[393];
assign   tb_i_rf_static_plaintext_length[394] =   64'h0000000000000280;
assign   tb_i_plaintext[394]                  =   tb_i_plaintext[393];
assign   tb_o_valid[394]                      =   1'b0;
assign   tb_o_sop[394]                        =   1'b0;
assign   tb_o_ciphertext[394]                 =   tb_o_ciphertext[393];
assign   tb_o_tag_ready[394]                  =   1'b0;
assign   tb_o_tag[394]                        =   tb_o_tag[393];

// CLK no. 395/1240
// *************************************************
assign   tb_i_valid[395]                      =   1'b0;
assign   tb_i_reset[395]                      =   1'b0;
assign   tb_i_sop[395]                        =   1'b0;
assign   tb_i_key_update[395]                 =   1'b0;
assign   tb_i_key[395]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[395]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[395]               =   1'b0;
assign   tb_i_rf_static_encrypt[395]          =   1'b1;
assign   tb_i_clear_fault_flags[395]          =   1'b0;
assign   tb_i_rf_static_aad_length[395]       =   64'h0000000000000100;
assign   tb_i_aad[395]                        =   tb_i_aad[394];
assign   tb_i_rf_static_plaintext_length[395] =   64'h0000000000000280;
assign   tb_i_plaintext[395]                  =   tb_i_plaintext[394];
assign   tb_o_valid[395]                      =   1'b0;
assign   tb_o_sop[395]                        =   1'b0;
assign   tb_o_ciphertext[395]                 =   tb_o_ciphertext[394];
assign   tb_o_tag_ready[395]                  =   1'b0;
assign   tb_o_tag[395]                        =   tb_o_tag[394];

// CLK no. 396/1240
// *************************************************
assign   tb_i_valid[396]                      =   1'b0;
assign   tb_i_reset[396]                      =   1'b0;
assign   tb_i_sop[396]                        =   1'b0;
assign   tb_i_key_update[396]                 =   1'b0;
assign   tb_i_key[396]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[396]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[396]               =   1'b0;
assign   tb_i_rf_static_encrypt[396]          =   1'b1;
assign   tb_i_clear_fault_flags[396]          =   1'b0;
assign   tb_i_rf_static_aad_length[396]       =   64'h0000000000000100;
assign   tb_i_aad[396]                        =   tb_i_aad[395];
assign   tb_i_rf_static_plaintext_length[396] =   64'h0000000000000280;
assign   tb_i_plaintext[396]                  =   tb_i_plaintext[395];
assign   tb_o_valid[396]                      =   1'b0;
assign   tb_o_sop[396]                        =   1'b0;
assign   tb_o_ciphertext[396]                 =   tb_o_ciphertext[395];
assign   tb_o_tag_ready[396]                  =   1'b0;
assign   tb_o_tag[396]                        =   tb_o_tag[395];

// CLK no. 397/1240
// *************************************************
assign   tb_i_valid[397]                      =   1'b0;
assign   tb_i_reset[397]                      =   1'b0;
assign   tb_i_sop[397]                        =   1'b0;
assign   tb_i_key_update[397]                 =   1'b0;
assign   tb_i_key[397]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[397]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[397]               =   1'b0;
assign   tb_i_rf_static_encrypt[397]          =   1'b1;
assign   tb_i_clear_fault_flags[397]          =   1'b0;
assign   tb_i_rf_static_aad_length[397]       =   64'h0000000000000100;
assign   tb_i_aad[397]                        =   tb_i_aad[396];
assign   tb_i_rf_static_plaintext_length[397] =   64'h0000000000000280;
assign   tb_i_plaintext[397]                  =   tb_i_plaintext[396];
assign   tb_o_valid[397]                      =   1'b0;
assign   tb_o_sop[397]                        =   1'b0;
assign   tb_o_ciphertext[397]                 =   tb_o_ciphertext[396];
assign   tb_o_tag_ready[397]                  =   1'b0;
assign   tb_o_tag[397]                        =   tb_o_tag[396];

// CLK no. 398/1240
// *************************************************
assign   tb_i_valid[398]                      =   1'b0;
assign   tb_i_reset[398]                      =   1'b0;
assign   tb_i_sop[398]                        =   1'b0;
assign   tb_i_key_update[398]                 =   1'b0;
assign   tb_i_key[398]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[398]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[398]               =   1'b0;
assign   tb_i_rf_static_encrypt[398]          =   1'b1;
assign   tb_i_clear_fault_flags[398]          =   1'b0;
assign   tb_i_rf_static_aad_length[398]       =   64'h0000000000000100;
assign   tb_i_aad[398]                        =   tb_i_aad[397];
assign   tb_i_rf_static_plaintext_length[398] =   64'h0000000000000280;
assign   tb_i_plaintext[398]                  =   tb_i_plaintext[397];
assign   tb_o_valid[398]                      =   1'b0;
assign   tb_o_sop[398]                        =   1'b0;
assign   tb_o_ciphertext[398]                 =   tb_o_ciphertext[397];
assign   tb_o_tag_ready[398]                  =   1'b0;
assign   tb_o_tag[398]                        =   tb_o_tag[397];

// CLK no. 399/1240
// *************************************************
assign   tb_i_valid[399]                      =   1'b0;
assign   tb_i_reset[399]                      =   1'b0;
assign   tb_i_sop[399]                        =   1'b0;
assign   tb_i_key_update[399]                 =   1'b0;
assign   tb_i_key[399]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[399]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[399]               =   1'b0;
assign   tb_i_rf_static_encrypt[399]          =   1'b1;
assign   tb_i_clear_fault_flags[399]          =   1'b0;
assign   tb_i_rf_static_aad_length[399]       =   64'h0000000000000100;
assign   tb_i_aad[399]                        =   tb_i_aad[398];
assign   tb_i_rf_static_plaintext_length[399] =   64'h0000000000000280;
assign   tb_i_plaintext[399]                  =   tb_i_plaintext[398];
assign   tb_o_valid[399]                      =   1'b0;
assign   tb_o_sop[399]                        =   1'b0;
assign   tb_o_ciphertext[399]                 =   tb_o_ciphertext[398];
assign   tb_o_tag_ready[399]                  =   1'b0;
assign   tb_o_tag[399]                        =   tb_o_tag[398];

// CLK no. 400/1240
// *************************************************
assign   tb_i_valid[400]                      =   1'b0;
assign   tb_i_reset[400]                      =   1'b0;
assign   tb_i_sop[400]                        =   1'b0;
assign   tb_i_key_update[400]                 =   1'b0;
assign   tb_i_key[400]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[400]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[400]               =   1'b0;
assign   tb_i_rf_static_encrypt[400]          =   1'b1;
assign   tb_i_clear_fault_flags[400]          =   1'b0;
assign   tb_i_rf_static_aad_length[400]       =   64'h0000000000000100;
assign   tb_i_aad[400]                        =   tb_i_aad[399];
assign   tb_i_rf_static_plaintext_length[400] =   64'h0000000000000280;
assign   tb_i_plaintext[400]                  =   tb_i_plaintext[399];
assign   tb_o_valid[400]                      =   1'b0;
assign   tb_o_sop[400]                        =   1'b0;
assign   tb_o_ciphertext[400]                 =   tb_o_ciphertext[399];
assign   tb_o_tag_ready[400]                  =   1'b0;
assign   tb_o_tag[400]                        =   tb_o_tag[399];

// CLK no. 401/1240
// *************************************************
assign   tb_i_valid[401]                      =   1'b0;
assign   tb_i_reset[401]                      =   1'b0;
assign   tb_i_sop[401]                        =   1'b0;
assign   tb_i_key_update[401]                 =   1'b0;
assign   tb_i_key[401]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[401]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[401]               =   1'b0;
assign   tb_i_rf_static_encrypt[401]          =   1'b1;
assign   tb_i_clear_fault_flags[401]          =   1'b0;
assign   tb_i_rf_static_aad_length[401]       =   64'h0000000000000100;
assign   tb_i_aad[401]                        =   tb_i_aad[400];
assign   tb_i_rf_static_plaintext_length[401] =   64'h0000000000000280;
assign   tb_i_plaintext[401]                  =   tb_i_plaintext[400];
assign   tb_o_valid[401]                      =   1'b1;
assign   tb_o_sop[401]                        =   1'b1;
assign   tb_o_ciphertext[401]                 =   256'hf4f842ee8b1b7b12778d6d3b807cd9ee5e6e264960002b5c16888a14af1a4581;
assign   tb_o_tag_ready[401]                  =   1'b0;
assign   tb_o_tag[401]                        =   tb_o_tag[400];

// CLK no. 402/1240
// *************************************************
assign   tb_i_valid[402]                      =   1'b0;
assign   tb_i_reset[402]                      =   1'b0;
assign   tb_i_sop[402]                        =   1'b0;
assign   tb_i_key_update[402]                 =   1'b0;
assign   tb_i_key[402]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[402]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[402]               =   1'b0;
assign   tb_i_rf_static_encrypt[402]          =   1'b1;
assign   tb_i_clear_fault_flags[402]          =   1'b0;
assign   tb_i_rf_static_aad_length[402]       =   64'h0000000000000100;
assign   tb_i_aad[402]                        =   tb_i_aad[401];
assign   tb_i_rf_static_plaintext_length[402] =   64'h0000000000000280;
assign   tb_i_plaintext[402]                  =   tb_i_plaintext[401];
assign   tb_o_valid[402]                      =   1'b1;
assign   tb_o_sop[402]                        =   1'b0;
assign   tb_o_ciphertext[402]                 =   256'hd965aa61d572756e75e8f5377c1eb112d028cebdb2b183c6e8dcf614087df7e0;
assign   tb_o_tag_ready[402]                  =   1'b0;
assign   tb_o_tag[402]                        =   tb_o_tag[401];

// CLK no. 403/1240
// *************************************************
assign   tb_i_valid[403]                      =   1'b0;
assign   tb_i_reset[403]                      =   1'b0;
assign   tb_i_sop[403]                        =   1'b0;
assign   tb_i_key_update[403]                 =   1'b0;
assign   tb_i_key[403]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[403]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[403]               =   1'b0;
assign   tb_i_rf_static_encrypt[403]          =   1'b1;
assign   tb_i_clear_fault_flags[403]          =   1'b0;
assign   tb_i_rf_static_aad_length[403]       =   64'h0000000000000100;
assign   tb_i_aad[403]                        =   tb_i_aad[402];
assign   tb_i_rf_static_plaintext_length[403] =   64'h0000000000000280;
assign   tb_i_plaintext[403]                  =   tb_i_plaintext[402];
assign   tb_o_valid[403]                      =   1'b1;
assign   tb_o_sop[403]                        =   1'b0;
assign   tb_o_ciphertext[403]                 =   256'had329d969b6850b333778804c56efb93;
assign   tb_o_tag_ready[403]                  =   1'b0;
assign   tb_o_tag[403]                        =   tb_o_tag[402];

// CLK no. 404/1240
// *************************************************
assign   tb_i_valid[404]                      =   1'b0;
assign   tb_i_reset[404]                      =   1'b0;
assign   tb_i_sop[404]                        =   1'b0;
assign   tb_i_key_update[404]                 =   1'b0;
assign   tb_i_key[404]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[404]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[404]               =   1'b0;
assign   tb_i_rf_static_encrypt[404]          =   1'b1;
assign   tb_i_clear_fault_flags[404]          =   1'b0;
assign   tb_i_rf_static_aad_length[404]       =   64'h0000000000000100;
assign   tb_i_aad[404]                        =   tb_i_aad[403];
assign   tb_i_rf_static_plaintext_length[404] =   64'h0000000000000280;
assign   tb_i_plaintext[404]                  =   tb_i_plaintext[403];
assign   tb_o_valid[404]                      =   1'b0;
assign   tb_o_sop[404]                        =   1'b0;
assign   tb_o_ciphertext[404]                 =   tb_o_ciphertext[403];
assign   tb_o_tag_ready[404]                  =   1'b0;
assign   tb_o_tag[404]                        =   tb_o_tag[403];

// CLK no. 405/1240
// *************************************************
assign   tb_i_valid[405]                      =   1'b0;
assign   tb_i_reset[405]                      =   1'b0;
assign   tb_i_sop[405]                        =   1'b0;
assign   tb_i_key_update[405]                 =   1'b0;
assign   tb_i_key[405]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[405]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[405]               =   1'b0;
assign   tb_i_rf_static_encrypt[405]          =   1'b1;
assign   tb_i_clear_fault_flags[405]          =   1'b0;
assign   tb_i_rf_static_aad_length[405]       =   64'h0000000000000100;
assign   tb_i_aad[405]                        =   tb_i_aad[404];
assign   tb_i_rf_static_plaintext_length[405] =   64'h0000000000000280;
assign   tb_i_plaintext[405]                  =   tb_i_plaintext[404];
assign   tb_o_valid[405]                      =   1'b0;
assign   tb_o_sop[405]                        =   1'b0;
assign   tb_o_ciphertext[405]                 =   tb_o_ciphertext[404];
assign   tb_o_tag_ready[405]                  =   1'b0;
assign   tb_o_tag[405]                        =   tb_o_tag[404];

// CLK no. 406/1240
// *************************************************
assign   tb_i_valid[406]                      =   1'b0;
assign   tb_i_reset[406]                      =   1'b0;
assign   tb_i_sop[406]                        =   1'b0;
assign   tb_i_key_update[406]                 =   1'b0;
assign   tb_i_key[406]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[406]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[406]               =   1'b0;
assign   tb_i_rf_static_encrypt[406]          =   1'b1;
assign   tb_i_clear_fault_flags[406]          =   1'b0;
assign   tb_i_rf_static_aad_length[406]       =   64'h0000000000000100;
assign   tb_i_aad[406]                        =   tb_i_aad[405];
assign   tb_i_rf_static_plaintext_length[406] =   64'h0000000000000280;
assign   tb_i_plaintext[406]                  =   tb_i_plaintext[405];
assign   tb_o_valid[406]                      =   1'b0;
assign   tb_o_sop[406]                        =   1'b0;
assign   tb_o_ciphertext[406]                 =   tb_o_ciphertext[405];
assign   tb_o_tag_ready[406]                  =   1'b0;
assign   tb_o_tag[406]                        =   tb_o_tag[405];

// CLK no. 407/1240
// *************************************************
assign   tb_i_valid[407]                      =   1'b0;
assign   tb_i_reset[407]                      =   1'b0;
assign   tb_i_sop[407]                        =   1'b0;
assign   tb_i_key_update[407]                 =   1'b0;
assign   tb_i_key[407]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[407]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[407]               =   1'b0;
assign   tb_i_rf_static_encrypt[407]          =   1'b1;
assign   tb_i_clear_fault_flags[407]          =   1'b0;
assign   tb_i_rf_static_aad_length[407]       =   64'h0000000000000100;
assign   tb_i_aad[407]                        =   tb_i_aad[406];
assign   tb_i_rf_static_plaintext_length[407] =   64'h0000000000000280;
assign   tb_i_plaintext[407]                  =   tb_i_plaintext[406];
assign   tb_o_valid[407]                      =   1'b0;
assign   tb_o_sop[407]                        =   1'b0;
assign   tb_o_ciphertext[407]                 =   tb_o_ciphertext[406];
assign   tb_o_tag_ready[407]                  =   1'b0;
assign   tb_o_tag[407]                        =   tb_o_tag[406];

// CLK no. 408/1240
// *************************************************
assign   tb_i_valid[408]                      =   1'b0;
assign   tb_i_reset[408]                      =   1'b0;
assign   tb_i_sop[408]                        =   1'b0;
assign   tb_i_key_update[408]                 =   1'b0;
assign   tb_i_key[408]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[408]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[408]               =   1'b0;
assign   tb_i_rf_static_encrypt[408]          =   1'b1;
assign   tb_i_clear_fault_flags[408]          =   1'b0;
assign   tb_i_rf_static_aad_length[408]       =   64'h0000000000000100;
assign   tb_i_aad[408]                        =   tb_i_aad[407];
assign   tb_i_rf_static_plaintext_length[408] =   64'h0000000000000280;
assign   tb_i_plaintext[408]                  =   tb_i_plaintext[407];
assign   tb_o_valid[408]                      =   1'b0;
assign   tb_o_sop[408]                        =   1'b0;
assign   tb_o_ciphertext[408]                 =   tb_o_ciphertext[407];
assign   tb_o_tag_ready[408]                  =   1'b0;
assign   tb_o_tag[408]                        =   tb_o_tag[407];

// CLK no. 409/1240
// *************************************************
assign   tb_i_valid[409]                      =   1'b0;
assign   tb_i_reset[409]                      =   1'b0;
assign   tb_i_sop[409]                        =   1'b0;
assign   tb_i_key_update[409]                 =   1'b0;
assign   tb_i_key[409]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[409]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[409]               =   1'b0;
assign   tb_i_rf_static_encrypt[409]          =   1'b1;
assign   tb_i_clear_fault_flags[409]          =   1'b0;
assign   tb_i_rf_static_aad_length[409]       =   64'h0000000000000100;
assign   tb_i_aad[409]                        =   tb_i_aad[408];
assign   tb_i_rf_static_plaintext_length[409] =   64'h0000000000000280;
assign   tb_i_plaintext[409]                  =   tb_i_plaintext[408];
assign   tb_o_valid[409]                      =   1'b0;
assign   tb_o_sop[409]                        =   1'b0;
assign   tb_o_ciphertext[409]                 =   tb_o_ciphertext[408];
assign   tb_o_tag_ready[409]                  =   1'b0;
assign   tb_o_tag[409]                        =   tb_o_tag[408];

// CLK no. 410/1240
// *************************************************
assign   tb_i_valid[410]                      =   1'b0;
assign   tb_i_reset[410]                      =   1'b0;
assign   tb_i_sop[410]                        =   1'b0;
assign   tb_i_key_update[410]                 =   1'b0;
assign   tb_i_key[410]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[410]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[410]               =   1'b0;
assign   tb_i_rf_static_encrypt[410]          =   1'b1;
assign   tb_i_clear_fault_flags[410]          =   1'b0;
assign   tb_i_rf_static_aad_length[410]       =   64'h0000000000000100;
assign   tb_i_aad[410]                        =   tb_i_aad[409];
assign   tb_i_rf_static_plaintext_length[410] =   64'h0000000000000280;
assign   tb_i_plaintext[410]                  =   tb_i_plaintext[409];
assign   tb_o_valid[410]                      =   1'b0;
assign   tb_o_sop[410]                        =   1'b0;
assign   tb_o_ciphertext[410]                 =   tb_o_ciphertext[409];
assign   tb_o_tag_ready[410]                  =   1'b0;
assign   tb_o_tag[410]                        =   tb_o_tag[409];

// CLK no. 411/1240
// *************************************************
assign   tb_i_valid[411]                      =   1'b0;
assign   tb_i_reset[411]                      =   1'b0;
assign   tb_i_sop[411]                        =   1'b0;
assign   tb_i_key_update[411]                 =   1'b0;
assign   tb_i_key[411]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[411]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[411]               =   1'b0;
assign   tb_i_rf_static_encrypt[411]          =   1'b1;
assign   tb_i_clear_fault_flags[411]          =   1'b0;
assign   tb_i_rf_static_aad_length[411]       =   64'h0000000000000100;
assign   tb_i_aad[411]                        =   tb_i_aad[410];
assign   tb_i_rf_static_plaintext_length[411] =   64'h0000000000000280;
assign   tb_i_plaintext[411]                  =   tb_i_plaintext[410];
assign   tb_o_valid[411]                      =   1'b0;
assign   tb_o_sop[411]                        =   1'b0;
assign   tb_o_ciphertext[411]                 =   tb_o_ciphertext[410];
assign   tb_o_tag_ready[411]                  =   1'b1;
assign   tb_o_tag[411]                        =   128'h1c4b5905b0c453050188b06ae6b7c2e7;

// CLK no. 412/1240
// *************************************************
assign   tb_i_valid[412]                      =   1'b0;
assign   tb_i_reset[412]                      =   1'b0;
assign   tb_i_sop[412]                        =   1'b0;
assign   tb_i_key_update[412]                 =   1'b0;
assign   tb_i_key[412]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[412]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[412]               =   1'b0;
assign   tb_i_rf_static_encrypt[412]          =   1'b1;
assign   tb_i_clear_fault_flags[412]          =   1'b0;
assign   tb_i_rf_static_aad_length[412]       =   64'h0000000000000100;
assign   tb_i_aad[412]                        =   tb_i_aad[411];
assign   tb_i_rf_static_plaintext_length[412] =   64'h0000000000000280;
assign   tb_i_plaintext[412]                  =   tb_i_plaintext[411];
assign   tb_o_valid[412]                      =   1'b0;
assign   tb_o_sop[412]                        =   1'b0;
assign   tb_o_ciphertext[412]                 =   tb_o_ciphertext[411];
assign   tb_o_tag_ready[412]                  =   1'b0;
assign   tb_o_tag[412]                        =   tb_o_tag[411];

// CLK no. 413/1240
// *************************************************
assign   tb_i_valid[413]                      =   1'b0;
assign   tb_i_reset[413]                      =   1'b0;
assign   tb_i_sop[413]                        =   1'b0;
assign   tb_i_key_update[413]                 =   1'b0;
assign   tb_i_key[413]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[413]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[413]               =   1'b0;
assign   tb_i_rf_static_encrypt[413]          =   1'b1;
assign   tb_i_clear_fault_flags[413]          =   1'b0;
assign   tb_i_rf_static_aad_length[413]       =   64'h0000000000000100;
assign   tb_i_aad[413]                        =   tb_i_aad[412];
assign   tb_i_rf_static_plaintext_length[413] =   64'h0000000000000280;
assign   tb_i_plaintext[413]                  =   tb_i_plaintext[412];
assign   tb_o_valid[413]                      =   1'b0;
assign   tb_o_sop[413]                        =   1'b0;
assign   tb_o_ciphertext[413]                 =   tb_o_ciphertext[412];
assign   tb_o_tag_ready[413]                  =   1'b0;
assign   tb_o_tag[413]                        =   tb_o_tag[412];

// CLK no. 414/1240
// *************************************************
assign   tb_i_valid[414]                      =   1'b0;
assign   tb_i_reset[414]                      =   1'b0;
assign   tb_i_sop[414]                        =   1'b1;
assign   tb_i_key_update[414]                 =   1'b0;
assign   tb_i_key[414]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[414]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[414]               =   1'b0;
assign   tb_i_rf_static_encrypt[414]          =   1'b1;
assign   tb_i_clear_fault_flags[414]          =   1'b0;
assign   tb_i_rf_static_aad_length[414]       =   64'h0000000000000100;
assign   tb_i_aad[414]                        =   tb_i_aad[413];
assign   tb_i_rf_static_plaintext_length[414] =   64'h0000000000000280;
assign   tb_i_plaintext[414]                  =   tb_i_plaintext[413];
assign   tb_o_valid[414]                      =   1'b0;
assign   tb_o_sop[414]                        =   1'b0;
assign   tb_o_ciphertext[414]                 =   tb_o_ciphertext[413];
assign   tb_o_tag_ready[414]                  =   1'b0;
assign   tb_o_tag[414]                        =   tb_o_tag[413];

// CLK no. 415/1240
// *************************************************
assign   tb_i_valid[415]                      =   1'b1;
assign   tb_i_reset[415]                      =   1'b0;
assign   tb_i_sop[415]                        =   1'b0;
assign   tb_i_key_update[415]                 =   1'b0;
assign   tb_i_key[415]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[415]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[415]               =   1'b0;
assign   tb_i_rf_static_encrypt[415]          =   1'b1;
assign   tb_i_clear_fault_flags[415]          =   1'b0;
assign   tb_i_rf_static_aad_length[415]       =   64'h0000000000000100;
assign   tb_i_aad[415]                        =   256'hd30c1db730e930a5fd26c518e5cf27b4248e79b5523ac09e693654c01b6c8147;
assign   tb_i_rf_static_plaintext_length[415] =   64'h0000000000000280;
assign   tb_i_plaintext[415]                  =   tb_i_plaintext[414];
assign   tb_o_valid[415]                      =   1'b0;
assign   tb_o_sop[415]                        =   1'b0;
assign   tb_o_ciphertext[415]                 =   tb_o_ciphertext[414];
assign   tb_o_tag_ready[415]                  =   1'b0;
assign   tb_o_tag[415]                        =   tb_o_tag[414];

// CLK no. 416/1240
// *************************************************
assign   tb_i_valid[416]                      =   1'b1;
assign   tb_i_reset[416]                      =   1'b0;
assign   tb_i_sop[416]                        =   1'b0;
assign   tb_i_key_update[416]                 =   1'b0;
assign   tb_i_key[416]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[416]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[416]               =   1'b0;
assign   tb_i_rf_static_encrypt[416]          =   1'b1;
assign   tb_i_clear_fault_flags[416]          =   1'b0;
assign   tb_i_rf_static_aad_length[416]       =   64'h0000000000000100;
assign   tb_i_aad[416]                        =   tb_i_aad[415];
assign   tb_i_rf_static_plaintext_length[416] =   64'h0000000000000280;
assign   tb_i_plaintext[416]                  =   256'h45899a688db97a2059ce9cfa0dd5bb29da16519d38cd1bc080c75ca26b82f997;
assign   tb_o_valid[416]                      =   1'b0;
assign   tb_o_sop[416]                        =   1'b0;
assign   tb_o_ciphertext[416]                 =   tb_o_ciphertext[415];
assign   tb_o_tag_ready[416]                  =   1'b0;
assign   tb_o_tag[416]                        =   tb_o_tag[415];

// CLK no. 417/1240
// *************************************************
assign   tb_i_valid[417]                      =   1'b1;
assign   tb_i_reset[417]                      =   1'b0;
assign   tb_i_sop[417]                        =   1'b0;
assign   tb_i_key_update[417]                 =   1'b0;
assign   tb_i_key[417]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[417]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[417]               =   1'b0;
assign   tb_i_rf_static_encrypt[417]          =   1'b1;
assign   tb_i_clear_fault_flags[417]          =   1'b0;
assign   tb_i_rf_static_aad_length[417]       =   64'h0000000000000100;
assign   tb_i_aad[417]                        =   tb_i_aad[416];
assign   tb_i_rf_static_plaintext_length[417] =   64'h0000000000000280;
assign   tb_i_plaintext[417]                  =   256'hd7f6f71304139687fa2e8556751d00c9f9611e8f38781149564ec456765d508b;
assign   tb_o_valid[417]                      =   1'b0;
assign   tb_o_sop[417]                        =   1'b0;
assign   tb_o_ciphertext[417]                 =   tb_o_ciphertext[416];
assign   tb_o_tag_ready[417]                  =   1'b0;
assign   tb_o_tag[417]                        =   tb_o_tag[416];

// CLK no. 418/1240
// *************************************************
assign   tb_i_valid[418]                      =   1'b1;
assign   tb_i_reset[418]                      =   1'b0;
assign   tb_i_sop[418]                        =   1'b0;
assign   tb_i_key_update[418]                 =   1'b0;
assign   tb_i_key[418]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[418]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[418]               =   1'b0;
assign   tb_i_rf_static_encrypt[418]          =   1'b1;
assign   tb_i_clear_fault_flags[418]          =   1'b0;
assign   tb_i_rf_static_aad_length[418]       =   64'h0000000000000100;
assign   tb_i_aad[418]                        =   tb_i_aad[417];
assign   tb_i_rf_static_plaintext_length[418] =   64'h0000000000000280;
assign   tb_i_plaintext[418]                  =   256'hc15891209d57adb6aae7b02cba2d0b8b;
assign   tb_o_valid[418]                      =   1'b0;
assign   tb_o_sop[418]                        =   1'b0;
assign   tb_o_ciphertext[418]                 =   tb_o_ciphertext[417];
assign   tb_o_tag_ready[418]                  =   1'b0;
assign   tb_o_tag[418]                        =   tb_o_tag[417];

// CLK no. 419/1240
// *************************************************
assign   tb_i_valid[419]                      =   1'b0;
assign   tb_i_reset[419]                      =   1'b0;
assign   tb_i_sop[419]                        =   1'b0;
assign   tb_i_key_update[419]                 =   1'b0;
assign   tb_i_key[419]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[419]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[419]               =   1'b0;
assign   tb_i_rf_static_encrypt[419]          =   1'b1;
assign   tb_i_clear_fault_flags[419]          =   1'b0;
assign   tb_i_rf_static_aad_length[419]       =   64'h0000000000000100;
assign   tb_i_aad[419]                        =   tb_i_aad[418];
assign   tb_i_rf_static_plaintext_length[419] =   64'h0000000000000280;
assign   tb_i_plaintext[419]                  =   tb_i_plaintext[418];
assign   tb_o_valid[419]                      =   1'b0;
assign   tb_o_sop[419]                        =   1'b0;
assign   tb_o_ciphertext[419]                 =   tb_o_ciphertext[418];
assign   tb_o_tag_ready[419]                  =   1'b0;
assign   tb_o_tag[419]                        =   tb_o_tag[418];

// CLK no. 420/1240
// *************************************************
assign   tb_i_valid[420]                      =   1'b0;
assign   tb_i_reset[420]                      =   1'b0;
assign   tb_i_sop[420]                        =   1'b0;
assign   tb_i_key_update[420]                 =   1'b0;
assign   tb_i_key[420]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[420]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[420]               =   1'b0;
assign   tb_i_rf_static_encrypt[420]          =   1'b1;
assign   tb_i_clear_fault_flags[420]          =   1'b0;
assign   tb_i_rf_static_aad_length[420]       =   64'h0000000000000100;
assign   tb_i_aad[420]                        =   tb_i_aad[419];
assign   tb_i_rf_static_plaintext_length[420] =   64'h0000000000000280;
assign   tb_i_plaintext[420]                  =   tb_i_plaintext[419];
assign   tb_o_valid[420]                      =   1'b0;
assign   tb_o_sop[420]                        =   1'b0;
assign   tb_o_ciphertext[420]                 =   tb_o_ciphertext[419];
assign   tb_o_tag_ready[420]                  =   1'b0;
assign   tb_o_tag[420]                        =   tb_o_tag[419];

// CLK no. 421/1240
// *************************************************
assign   tb_i_valid[421]                      =   1'b0;
assign   tb_i_reset[421]                      =   1'b0;
assign   tb_i_sop[421]                        =   1'b0;
assign   tb_i_key_update[421]                 =   1'b0;
assign   tb_i_key[421]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[421]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[421]               =   1'b0;
assign   tb_i_rf_static_encrypt[421]          =   1'b1;
assign   tb_i_clear_fault_flags[421]          =   1'b0;
assign   tb_i_rf_static_aad_length[421]       =   64'h0000000000000100;
assign   tb_i_aad[421]                        =   tb_i_aad[420];
assign   tb_i_rf_static_plaintext_length[421] =   64'h0000000000000280;
assign   tb_i_plaintext[421]                  =   tb_i_plaintext[420];
assign   tb_o_valid[421]                      =   1'b0;
assign   tb_o_sop[421]                        =   1'b0;
assign   tb_o_ciphertext[421]                 =   tb_o_ciphertext[420];
assign   tb_o_tag_ready[421]                  =   1'b0;
assign   tb_o_tag[421]                        =   tb_o_tag[420];

// CLK no. 422/1240
// *************************************************
assign   tb_i_valid[422]                      =   1'b0;
assign   tb_i_reset[422]                      =   1'b0;
assign   tb_i_sop[422]                        =   1'b0;
assign   tb_i_key_update[422]                 =   1'b0;
assign   tb_i_key[422]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[422]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[422]               =   1'b0;
assign   tb_i_rf_static_encrypt[422]          =   1'b1;
assign   tb_i_clear_fault_flags[422]          =   1'b0;
assign   tb_i_rf_static_aad_length[422]       =   64'h0000000000000100;
assign   tb_i_aad[422]                        =   tb_i_aad[421];
assign   tb_i_rf_static_plaintext_length[422] =   64'h0000000000000280;
assign   tb_i_plaintext[422]                  =   tb_i_plaintext[421];
assign   tb_o_valid[422]                      =   1'b0;
assign   tb_o_sop[422]                        =   1'b0;
assign   tb_o_ciphertext[422]                 =   tb_o_ciphertext[421];
assign   tb_o_tag_ready[422]                  =   1'b0;
assign   tb_o_tag[422]                        =   tb_o_tag[421];

// CLK no. 423/1240
// *************************************************
assign   tb_i_valid[423]                      =   1'b0;
assign   tb_i_reset[423]                      =   1'b0;
assign   tb_i_sop[423]                        =   1'b0;
assign   tb_i_key_update[423]                 =   1'b0;
assign   tb_i_key[423]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[423]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[423]               =   1'b0;
assign   tb_i_rf_static_encrypt[423]          =   1'b1;
assign   tb_i_clear_fault_flags[423]          =   1'b0;
assign   tb_i_rf_static_aad_length[423]       =   64'h0000000000000100;
assign   tb_i_aad[423]                        =   tb_i_aad[422];
assign   tb_i_rf_static_plaintext_length[423] =   64'h0000000000000280;
assign   tb_i_plaintext[423]                  =   tb_i_plaintext[422];
assign   tb_o_valid[423]                      =   1'b0;
assign   tb_o_sop[423]                        =   1'b0;
assign   tb_o_ciphertext[423]                 =   tb_o_ciphertext[422];
assign   tb_o_tag_ready[423]                  =   1'b0;
assign   tb_o_tag[423]                        =   tb_o_tag[422];

// CLK no. 424/1240
// *************************************************
assign   tb_i_valid[424]                      =   1'b0;
assign   tb_i_reset[424]                      =   1'b0;
assign   tb_i_sop[424]                        =   1'b0;
assign   tb_i_key_update[424]                 =   1'b0;
assign   tb_i_key[424]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[424]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[424]               =   1'b0;
assign   tb_i_rf_static_encrypt[424]          =   1'b1;
assign   tb_i_clear_fault_flags[424]          =   1'b0;
assign   tb_i_rf_static_aad_length[424]       =   64'h0000000000000100;
assign   tb_i_aad[424]                        =   tb_i_aad[423];
assign   tb_i_rf_static_plaintext_length[424] =   64'h0000000000000280;
assign   tb_i_plaintext[424]                  =   tb_i_plaintext[423];
assign   tb_o_valid[424]                      =   1'b0;
assign   tb_o_sop[424]                        =   1'b0;
assign   tb_o_ciphertext[424]                 =   tb_o_ciphertext[423];
assign   tb_o_tag_ready[424]                  =   1'b0;
assign   tb_o_tag[424]                        =   tb_o_tag[423];

// CLK no. 425/1240
// *************************************************
assign   tb_i_valid[425]                      =   1'b0;
assign   tb_i_reset[425]                      =   1'b0;
assign   tb_i_sop[425]                        =   1'b0;
assign   tb_i_key_update[425]                 =   1'b0;
assign   tb_i_key[425]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[425]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[425]               =   1'b0;
assign   tb_i_rf_static_encrypt[425]          =   1'b1;
assign   tb_i_clear_fault_flags[425]          =   1'b0;
assign   tb_i_rf_static_aad_length[425]       =   64'h0000000000000100;
assign   tb_i_aad[425]                        =   tb_i_aad[424];
assign   tb_i_rf_static_plaintext_length[425] =   64'h0000000000000280;
assign   tb_i_plaintext[425]                  =   tb_i_plaintext[424];
assign   tb_o_valid[425]                      =   1'b0;
assign   tb_o_sop[425]                        =   1'b0;
assign   tb_o_ciphertext[425]                 =   tb_o_ciphertext[424];
assign   tb_o_tag_ready[425]                  =   1'b0;
assign   tb_o_tag[425]                        =   tb_o_tag[424];

// CLK no. 426/1240
// *************************************************
assign   tb_i_valid[426]                      =   1'b0;
assign   tb_i_reset[426]                      =   1'b0;
assign   tb_i_sop[426]                        =   1'b0;
assign   tb_i_key_update[426]                 =   1'b0;
assign   tb_i_key[426]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[426]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[426]               =   1'b0;
assign   tb_i_rf_static_encrypt[426]          =   1'b1;
assign   tb_i_clear_fault_flags[426]          =   1'b0;
assign   tb_i_rf_static_aad_length[426]       =   64'h0000000000000100;
assign   tb_i_aad[426]                        =   tb_i_aad[425];
assign   tb_i_rf_static_plaintext_length[426] =   64'h0000000000000280;
assign   tb_i_plaintext[426]                  =   tb_i_plaintext[425];
assign   tb_o_valid[426]                      =   1'b0;
assign   tb_o_sop[426]                        =   1'b0;
assign   tb_o_ciphertext[426]                 =   tb_o_ciphertext[425];
assign   tb_o_tag_ready[426]                  =   1'b0;
assign   tb_o_tag[426]                        =   tb_o_tag[425];

// CLK no. 427/1240
// *************************************************
assign   tb_i_valid[427]                      =   1'b0;
assign   tb_i_reset[427]                      =   1'b0;
assign   tb_i_sop[427]                        =   1'b0;
assign   tb_i_key_update[427]                 =   1'b0;
assign   tb_i_key[427]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[427]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[427]               =   1'b0;
assign   tb_i_rf_static_encrypt[427]          =   1'b1;
assign   tb_i_clear_fault_flags[427]          =   1'b0;
assign   tb_i_rf_static_aad_length[427]       =   64'h0000000000000100;
assign   tb_i_aad[427]                        =   tb_i_aad[426];
assign   tb_i_rf_static_plaintext_length[427] =   64'h0000000000000280;
assign   tb_i_plaintext[427]                  =   tb_i_plaintext[426];
assign   tb_o_valid[427]                      =   1'b0;
assign   tb_o_sop[427]                        =   1'b0;
assign   tb_o_ciphertext[427]                 =   tb_o_ciphertext[426];
assign   tb_o_tag_ready[427]                  =   1'b0;
assign   tb_o_tag[427]                        =   tb_o_tag[426];

// CLK no. 428/1240
// *************************************************
assign   tb_i_valid[428]                      =   1'b0;
assign   tb_i_reset[428]                      =   1'b0;
assign   tb_i_sop[428]                        =   1'b0;
assign   tb_i_key_update[428]                 =   1'b0;
assign   tb_i_key[428]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[428]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[428]               =   1'b0;
assign   tb_i_rf_static_encrypt[428]          =   1'b1;
assign   tb_i_clear_fault_flags[428]          =   1'b0;
assign   tb_i_rf_static_aad_length[428]       =   64'h0000000000000100;
assign   tb_i_aad[428]                        =   tb_i_aad[427];
assign   tb_i_rf_static_plaintext_length[428] =   64'h0000000000000280;
assign   tb_i_plaintext[428]                  =   tb_i_plaintext[427];
assign   tb_o_valid[428]                      =   1'b0;
assign   tb_o_sop[428]                        =   1'b0;
assign   tb_o_ciphertext[428]                 =   tb_o_ciphertext[427];
assign   tb_o_tag_ready[428]                  =   1'b0;
assign   tb_o_tag[428]                        =   tb_o_tag[427];

// CLK no. 429/1240
// *************************************************
assign   tb_i_valid[429]                      =   1'b0;
assign   tb_i_reset[429]                      =   1'b0;
assign   tb_i_sop[429]                        =   1'b0;
assign   tb_i_key_update[429]                 =   1'b0;
assign   tb_i_key[429]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[429]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[429]               =   1'b0;
assign   tb_i_rf_static_encrypt[429]          =   1'b1;
assign   tb_i_clear_fault_flags[429]          =   1'b0;
assign   tb_i_rf_static_aad_length[429]       =   64'h0000000000000100;
assign   tb_i_aad[429]                        =   tb_i_aad[428];
assign   tb_i_rf_static_plaintext_length[429] =   64'h0000000000000280;
assign   tb_i_plaintext[429]                  =   tb_i_plaintext[428];
assign   tb_o_valid[429]                      =   1'b0;
assign   tb_o_sop[429]                        =   1'b0;
assign   tb_o_ciphertext[429]                 =   tb_o_ciphertext[428];
assign   tb_o_tag_ready[429]                  =   1'b0;
assign   tb_o_tag[429]                        =   tb_o_tag[428];

// CLK no. 430/1240
// *************************************************
assign   tb_i_valid[430]                      =   1'b0;
assign   tb_i_reset[430]                      =   1'b0;
assign   tb_i_sop[430]                        =   1'b0;
assign   tb_i_key_update[430]                 =   1'b0;
assign   tb_i_key[430]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[430]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[430]               =   1'b0;
assign   tb_i_rf_static_encrypt[430]          =   1'b1;
assign   tb_i_clear_fault_flags[430]          =   1'b0;
assign   tb_i_rf_static_aad_length[430]       =   64'h0000000000000100;
assign   tb_i_aad[430]                        =   tb_i_aad[429];
assign   tb_i_rf_static_plaintext_length[430] =   64'h0000000000000280;
assign   tb_i_plaintext[430]                  =   tb_i_plaintext[429];
assign   tb_o_valid[430]                      =   1'b0;
assign   tb_o_sop[430]                        =   1'b0;
assign   tb_o_ciphertext[430]                 =   tb_o_ciphertext[429];
assign   tb_o_tag_ready[430]                  =   1'b0;
assign   tb_o_tag[430]                        =   tb_o_tag[429];

// CLK no. 431/1240
// *************************************************
assign   tb_i_valid[431]                      =   1'b0;
assign   tb_i_reset[431]                      =   1'b0;
assign   tb_i_sop[431]                        =   1'b0;
assign   tb_i_key_update[431]                 =   1'b0;
assign   tb_i_key[431]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[431]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[431]               =   1'b0;
assign   tb_i_rf_static_encrypt[431]          =   1'b1;
assign   tb_i_clear_fault_flags[431]          =   1'b0;
assign   tb_i_rf_static_aad_length[431]       =   64'h0000000000000100;
assign   tb_i_aad[431]                        =   tb_i_aad[430];
assign   tb_i_rf_static_plaintext_length[431] =   64'h0000000000000280;
assign   tb_i_plaintext[431]                  =   tb_i_plaintext[430];
assign   tb_o_valid[431]                      =   1'b0;
assign   tb_o_sop[431]                        =   1'b0;
assign   tb_o_ciphertext[431]                 =   tb_o_ciphertext[430];
assign   tb_o_tag_ready[431]                  =   1'b0;
assign   tb_o_tag[431]                        =   tb_o_tag[430];

// CLK no. 432/1240
// *************************************************
assign   tb_i_valid[432]                      =   1'b0;
assign   tb_i_reset[432]                      =   1'b0;
assign   tb_i_sop[432]                        =   1'b0;
assign   tb_i_key_update[432]                 =   1'b0;
assign   tb_i_key[432]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[432]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[432]               =   1'b0;
assign   tb_i_rf_static_encrypt[432]          =   1'b1;
assign   tb_i_clear_fault_flags[432]          =   1'b0;
assign   tb_i_rf_static_aad_length[432]       =   64'h0000000000000100;
assign   tb_i_aad[432]                        =   tb_i_aad[431];
assign   tb_i_rf_static_plaintext_length[432] =   64'h0000000000000280;
assign   tb_i_plaintext[432]                  =   tb_i_plaintext[431];
assign   tb_o_valid[432]                      =   1'b0;
assign   tb_o_sop[432]                        =   1'b0;
assign   tb_o_ciphertext[432]                 =   tb_o_ciphertext[431];
assign   tb_o_tag_ready[432]                  =   1'b0;
assign   tb_o_tag[432]                        =   tb_o_tag[431];

// CLK no. 433/1240
// *************************************************
assign   tb_i_valid[433]                      =   1'b0;
assign   tb_i_reset[433]                      =   1'b0;
assign   tb_i_sop[433]                        =   1'b0;
assign   tb_i_key_update[433]                 =   1'b0;
assign   tb_i_key[433]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[433]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[433]               =   1'b0;
assign   tb_i_rf_static_encrypt[433]          =   1'b1;
assign   tb_i_clear_fault_flags[433]          =   1'b0;
assign   tb_i_rf_static_aad_length[433]       =   64'h0000000000000100;
assign   tb_i_aad[433]                        =   tb_i_aad[432];
assign   tb_i_rf_static_plaintext_length[433] =   64'h0000000000000280;
assign   tb_i_plaintext[433]                  =   tb_i_plaintext[432];
assign   tb_o_valid[433]                      =   1'b0;
assign   tb_o_sop[433]                        =   1'b0;
assign   tb_o_ciphertext[433]                 =   tb_o_ciphertext[432];
assign   tb_o_tag_ready[433]                  =   1'b0;
assign   tb_o_tag[433]                        =   tb_o_tag[432];

// CLK no. 434/1240
// *************************************************
assign   tb_i_valid[434]                      =   1'b0;
assign   tb_i_reset[434]                      =   1'b0;
assign   tb_i_sop[434]                        =   1'b0;
assign   tb_i_key_update[434]                 =   1'b0;
assign   tb_i_key[434]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[434]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[434]               =   1'b0;
assign   tb_i_rf_static_encrypt[434]          =   1'b1;
assign   tb_i_clear_fault_flags[434]          =   1'b0;
assign   tb_i_rf_static_aad_length[434]       =   64'h0000000000000100;
assign   tb_i_aad[434]                        =   tb_i_aad[433];
assign   tb_i_rf_static_plaintext_length[434] =   64'h0000000000000280;
assign   tb_i_plaintext[434]                  =   tb_i_plaintext[433];
assign   tb_o_valid[434]                      =   1'b0;
assign   tb_o_sop[434]                        =   1'b0;
assign   tb_o_ciphertext[434]                 =   tb_o_ciphertext[433];
assign   tb_o_tag_ready[434]                  =   1'b0;
assign   tb_o_tag[434]                        =   tb_o_tag[433];

// CLK no. 435/1240
// *************************************************
assign   tb_i_valid[435]                      =   1'b0;
assign   tb_i_reset[435]                      =   1'b0;
assign   tb_i_sop[435]                        =   1'b0;
assign   tb_i_key_update[435]                 =   1'b0;
assign   tb_i_key[435]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[435]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[435]               =   1'b0;
assign   tb_i_rf_static_encrypt[435]          =   1'b1;
assign   tb_i_clear_fault_flags[435]          =   1'b0;
assign   tb_i_rf_static_aad_length[435]       =   64'h0000000000000100;
assign   tb_i_aad[435]                        =   tb_i_aad[434];
assign   tb_i_rf_static_plaintext_length[435] =   64'h0000000000000280;
assign   tb_i_plaintext[435]                  =   tb_i_plaintext[434];
assign   tb_o_valid[435]                      =   1'b0;
assign   tb_o_sop[435]                        =   1'b0;
assign   tb_o_ciphertext[435]                 =   tb_o_ciphertext[434];
assign   tb_o_tag_ready[435]                  =   1'b0;
assign   tb_o_tag[435]                        =   tb_o_tag[434];

// CLK no. 436/1240
// *************************************************
assign   tb_i_valid[436]                      =   1'b0;
assign   tb_i_reset[436]                      =   1'b0;
assign   tb_i_sop[436]                        =   1'b0;
assign   tb_i_key_update[436]                 =   1'b0;
assign   tb_i_key[436]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[436]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[436]               =   1'b0;
assign   tb_i_rf_static_encrypt[436]          =   1'b1;
assign   tb_i_clear_fault_flags[436]          =   1'b0;
assign   tb_i_rf_static_aad_length[436]       =   64'h0000000000000100;
assign   tb_i_aad[436]                        =   tb_i_aad[435];
assign   tb_i_rf_static_plaintext_length[436] =   64'h0000000000000280;
assign   tb_i_plaintext[436]                  =   tb_i_plaintext[435];
assign   tb_o_valid[436]                      =   1'b0;
assign   tb_o_sop[436]                        =   1'b0;
assign   tb_o_ciphertext[436]                 =   tb_o_ciphertext[435];
assign   tb_o_tag_ready[436]                  =   1'b0;
assign   tb_o_tag[436]                        =   tb_o_tag[435];

// CLK no. 437/1240
// *************************************************
assign   tb_i_valid[437]                      =   1'b0;
assign   tb_i_reset[437]                      =   1'b0;
assign   tb_i_sop[437]                        =   1'b0;
assign   tb_i_key_update[437]                 =   1'b0;
assign   tb_i_key[437]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[437]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[437]               =   1'b0;
assign   tb_i_rf_static_encrypt[437]          =   1'b1;
assign   tb_i_clear_fault_flags[437]          =   1'b0;
assign   tb_i_rf_static_aad_length[437]       =   64'h0000000000000100;
assign   tb_i_aad[437]                        =   tb_i_aad[436];
assign   tb_i_rf_static_plaintext_length[437] =   64'h0000000000000280;
assign   tb_i_plaintext[437]                  =   tb_i_plaintext[436];
assign   tb_o_valid[437]                      =   1'b0;
assign   tb_o_sop[437]                        =   1'b0;
assign   tb_o_ciphertext[437]                 =   tb_o_ciphertext[436];
assign   tb_o_tag_ready[437]                  =   1'b0;
assign   tb_o_tag[437]                        =   tb_o_tag[436];

// CLK no. 438/1240
// *************************************************
assign   tb_i_valid[438]                      =   1'b0;
assign   tb_i_reset[438]                      =   1'b0;
assign   tb_i_sop[438]                        =   1'b0;
assign   tb_i_key_update[438]                 =   1'b0;
assign   tb_i_key[438]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[438]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[438]               =   1'b0;
assign   tb_i_rf_static_encrypt[438]          =   1'b1;
assign   tb_i_clear_fault_flags[438]          =   1'b0;
assign   tb_i_rf_static_aad_length[438]       =   64'h0000000000000100;
assign   tb_i_aad[438]                        =   tb_i_aad[437];
assign   tb_i_rf_static_plaintext_length[438] =   64'h0000000000000280;
assign   tb_i_plaintext[438]                  =   tb_i_plaintext[437];
assign   tb_o_valid[438]                      =   1'b0;
assign   tb_o_sop[438]                        =   1'b0;
assign   tb_o_ciphertext[438]                 =   tb_o_ciphertext[437];
assign   tb_o_tag_ready[438]                  =   1'b0;
assign   tb_o_tag[438]                        =   tb_o_tag[437];

// CLK no. 439/1240
// *************************************************
assign   tb_i_valid[439]                      =   1'b0;
assign   tb_i_reset[439]                      =   1'b0;
assign   tb_i_sop[439]                        =   1'b0;
assign   tb_i_key_update[439]                 =   1'b0;
assign   tb_i_key[439]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[439]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[439]               =   1'b0;
assign   tb_i_rf_static_encrypt[439]          =   1'b1;
assign   tb_i_clear_fault_flags[439]          =   1'b0;
assign   tb_i_rf_static_aad_length[439]       =   64'h0000000000000100;
assign   tb_i_aad[439]                        =   tb_i_aad[438];
assign   tb_i_rf_static_plaintext_length[439] =   64'h0000000000000280;
assign   tb_i_plaintext[439]                  =   tb_i_plaintext[438];
assign   tb_o_valid[439]                      =   1'b0;
assign   tb_o_sop[439]                        =   1'b0;
assign   tb_o_ciphertext[439]                 =   tb_o_ciphertext[438];
assign   tb_o_tag_ready[439]                  =   1'b0;
assign   tb_o_tag[439]                        =   tb_o_tag[438];

// CLK no. 440/1240
// *************************************************
assign   tb_i_valid[440]                      =   1'b0;
assign   tb_i_reset[440]                      =   1'b0;
assign   tb_i_sop[440]                        =   1'b0;
assign   tb_i_key_update[440]                 =   1'b0;
assign   tb_i_key[440]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[440]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[440]               =   1'b0;
assign   tb_i_rf_static_encrypt[440]          =   1'b1;
assign   tb_i_clear_fault_flags[440]          =   1'b0;
assign   tb_i_rf_static_aad_length[440]       =   64'h0000000000000100;
assign   tb_i_aad[440]                        =   tb_i_aad[439];
assign   tb_i_rf_static_plaintext_length[440] =   64'h0000000000000280;
assign   tb_i_plaintext[440]                  =   tb_i_plaintext[439];
assign   tb_o_valid[440]                      =   1'b0;
assign   tb_o_sop[440]                        =   1'b0;
assign   tb_o_ciphertext[440]                 =   tb_o_ciphertext[439];
assign   tb_o_tag_ready[440]                  =   1'b0;
assign   tb_o_tag[440]                        =   tb_o_tag[439];

// CLK no. 441/1240
// *************************************************
assign   tb_i_valid[441]                      =   1'b0;
assign   tb_i_reset[441]                      =   1'b0;
assign   tb_i_sop[441]                        =   1'b0;
assign   tb_i_key_update[441]                 =   1'b0;
assign   tb_i_key[441]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[441]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[441]               =   1'b0;
assign   tb_i_rf_static_encrypt[441]          =   1'b1;
assign   tb_i_clear_fault_flags[441]          =   1'b0;
assign   tb_i_rf_static_aad_length[441]       =   64'h0000000000000100;
assign   tb_i_aad[441]                        =   tb_i_aad[440];
assign   tb_i_rf_static_plaintext_length[441] =   64'h0000000000000280;
assign   tb_i_plaintext[441]                  =   tb_i_plaintext[440];
assign   tb_o_valid[441]                      =   1'b0;
assign   tb_o_sop[441]                        =   1'b0;
assign   tb_o_ciphertext[441]                 =   tb_o_ciphertext[440];
assign   tb_o_tag_ready[441]                  =   1'b0;
assign   tb_o_tag[441]                        =   tb_o_tag[440];

// CLK no. 442/1240
// *************************************************
assign   tb_i_valid[442]                      =   1'b0;
assign   tb_i_reset[442]                      =   1'b0;
assign   tb_i_sop[442]                        =   1'b0;
assign   tb_i_key_update[442]                 =   1'b0;
assign   tb_i_key[442]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[442]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[442]               =   1'b0;
assign   tb_i_rf_static_encrypt[442]          =   1'b1;
assign   tb_i_clear_fault_flags[442]          =   1'b0;
assign   tb_i_rf_static_aad_length[442]       =   64'h0000000000000100;
assign   tb_i_aad[442]                        =   tb_i_aad[441];
assign   tb_i_rf_static_plaintext_length[442] =   64'h0000000000000280;
assign   tb_i_plaintext[442]                  =   tb_i_plaintext[441];
assign   tb_o_valid[442]                      =   1'b0;
assign   tb_o_sop[442]                        =   1'b0;
assign   tb_o_ciphertext[442]                 =   tb_o_ciphertext[441];
assign   tb_o_tag_ready[442]                  =   1'b0;
assign   tb_o_tag[442]                        =   tb_o_tag[441];

// CLK no. 443/1240
// *************************************************
assign   tb_i_valid[443]                      =   1'b0;
assign   tb_i_reset[443]                      =   1'b0;
assign   tb_i_sop[443]                        =   1'b0;
assign   tb_i_key_update[443]                 =   1'b0;
assign   tb_i_key[443]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[443]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[443]               =   1'b0;
assign   tb_i_rf_static_encrypt[443]          =   1'b1;
assign   tb_i_clear_fault_flags[443]          =   1'b0;
assign   tb_i_rf_static_aad_length[443]       =   64'h0000000000000100;
assign   tb_i_aad[443]                        =   tb_i_aad[442];
assign   tb_i_rf_static_plaintext_length[443] =   64'h0000000000000280;
assign   tb_i_plaintext[443]                  =   tb_i_plaintext[442];
assign   tb_o_valid[443]                      =   1'b0;
assign   tb_o_sop[443]                        =   1'b0;
assign   tb_o_ciphertext[443]                 =   tb_o_ciphertext[442];
assign   tb_o_tag_ready[443]                  =   1'b0;
assign   tb_o_tag[443]                        =   tb_o_tag[442];

// CLK no. 444/1240
// *************************************************
assign   tb_i_valid[444]                      =   1'b0;
assign   tb_i_reset[444]                      =   1'b0;
assign   tb_i_sop[444]                        =   1'b0;
assign   tb_i_key_update[444]                 =   1'b0;
assign   tb_i_key[444]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[444]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[444]               =   1'b0;
assign   tb_i_rf_static_encrypt[444]          =   1'b1;
assign   tb_i_clear_fault_flags[444]          =   1'b0;
assign   tb_i_rf_static_aad_length[444]       =   64'h0000000000000100;
assign   tb_i_aad[444]                        =   tb_i_aad[443];
assign   tb_i_rf_static_plaintext_length[444] =   64'h0000000000000280;
assign   tb_i_plaintext[444]                  =   tb_i_plaintext[443];
assign   tb_o_valid[444]                      =   1'b0;
assign   tb_o_sop[444]                        =   1'b0;
assign   tb_o_ciphertext[444]                 =   tb_o_ciphertext[443];
assign   tb_o_tag_ready[444]                  =   1'b0;
assign   tb_o_tag[444]                        =   tb_o_tag[443];

// CLK no. 445/1240
// *************************************************
assign   tb_i_valid[445]                      =   1'b0;
assign   tb_i_reset[445]                      =   1'b0;
assign   tb_i_sop[445]                        =   1'b0;
assign   tb_i_key_update[445]                 =   1'b0;
assign   tb_i_key[445]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[445]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[445]               =   1'b0;
assign   tb_i_rf_static_encrypt[445]          =   1'b1;
assign   tb_i_clear_fault_flags[445]          =   1'b0;
assign   tb_i_rf_static_aad_length[445]       =   64'h0000000000000100;
assign   tb_i_aad[445]                        =   tb_i_aad[444];
assign   tb_i_rf_static_plaintext_length[445] =   64'h0000000000000280;
assign   tb_i_plaintext[445]                  =   tb_i_plaintext[444];
assign   tb_o_valid[445]                      =   1'b0;
assign   tb_o_sop[445]                        =   1'b0;
assign   tb_o_ciphertext[445]                 =   tb_o_ciphertext[444];
assign   tb_o_tag_ready[445]                  =   1'b0;
assign   tb_o_tag[445]                        =   tb_o_tag[444];

// CLK no. 446/1240
// *************************************************
assign   tb_i_valid[446]                      =   1'b0;
assign   tb_i_reset[446]                      =   1'b0;
assign   tb_i_sop[446]                        =   1'b0;
assign   tb_i_key_update[446]                 =   1'b0;
assign   tb_i_key[446]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[446]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[446]               =   1'b0;
assign   tb_i_rf_static_encrypt[446]          =   1'b1;
assign   tb_i_clear_fault_flags[446]          =   1'b0;
assign   tb_i_rf_static_aad_length[446]       =   64'h0000000000000100;
assign   tb_i_aad[446]                        =   tb_i_aad[445];
assign   tb_i_rf_static_plaintext_length[446] =   64'h0000000000000280;
assign   tb_i_plaintext[446]                  =   tb_i_plaintext[445];
assign   tb_o_valid[446]                      =   1'b0;
assign   tb_o_sop[446]                        =   1'b0;
assign   tb_o_ciphertext[446]                 =   tb_o_ciphertext[445];
assign   tb_o_tag_ready[446]                  =   1'b0;
assign   tb_o_tag[446]                        =   tb_o_tag[445];

// CLK no. 447/1240
// *************************************************
assign   tb_i_valid[447]                      =   1'b0;
assign   tb_i_reset[447]                      =   1'b0;
assign   tb_i_sop[447]                        =   1'b0;
assign   tb_i_key_update[447]                 =   1'b0;
assign   tb_i_key[447]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[447]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[447]               =   1'b0;
assign   tb_i_rf_static_encrypt[447]          =   1'b1;
assign   tb_i_clear_fault_flags[447]          =   1'b0;
assign   tb_i_rf_static_aad_length[447]       =   64'h0000000000000100;
assign   tb_i_aad[447]                        =   tb_i_aad[446];
assign   tb_i_rf_static_plaintext_length[447] =   64'h0000000000000280;
assign   tb_i_plaintext[447]                  =   tb_i_plaintext[446];
assign   tb_o_valid[447]                      =   1'b0;
assign   tb_o_sop[447]                        =   1'b0;
assign   tb_o_ciphertext[447]                 =   tb_o_ciphertext[446];
assign   tb_o_tag_ready[447]                  =   1'b0;
assign   tb_o_tag[447]                        =   tb_o_tag[446];

// CLK no. 448/1240
// *************************************************
assign   tb_i_valid[448]                      =   1'b0;
assign   tb_i_reset[448]                      =   1'b0;
assign   tb_i_sop[448]                        =   1'b0;
assign   tb_i_key_update[448]                 =   1'b0;
assign   tb_i_key[448]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[448]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[448]               =   1'b0;
assign   tb_i_rf_static_encrypt[448]          =   1'b1;
assign   tb_i_clear_fault_flags[448]          =   1'b0;
assign   tb_i_rf_static_aad_length[448]       =   64'h0000000000000100;
assign   tb_i_aad[448]                        =   tb_i_aad[447];
assign   tb_i_rf_static_plaintext_length[448] =   64'h0000000000000280;
assign   tb_i_plaintext[448]                  =   tb_i_plaintext[447];
assign   tb_o_valid[448]                      =   1'b0;
assign   tb_o_sop[448]                        =   1'b0;
assign   tb_o_ciphertext[448]                 =   tb_o_ciphertext[447];
assign   tb_o_tag_ready[448]                  =   1'b0;
assign   tb_o_tag[448]                        =   tb_o_tag[447];

// CLK no. 449/1240
// *************************************************
assign   tb_i_valid[449]                      =   1'b0;
assign   tb_i_reset[449]                      =   1'b0;
assign   tb_i_sop[449]                        =   1'b0;
assign   tb_i_key_update[449]                 =   1'b0;
assign   tb_i_key[449]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[449]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[449]               =   1'b0;
assign   tb_i_rf_static_encrypt[449]          =   1'b1;
assign   tb_i_clear_fault_flags[449]          =   1'b0;
assign   tb_i_rf_static_aad_length[449]       =   64'h0000000000000100;
assign   tb_i_aad[449]                        =   tb_i_aad[448];
assign   tb_i_rf_static_plaintext_length[449] =   64'h0000000000000280;
assign   tb_i_plaintext[449]                  =   tb_i_plaintext[448];
assign   tb_o_valid[449]                      =   1'b0;
assign   tb_o_sop[449]                        =   1'b0;
assign   tb_o_ciphertext[449]                 =   tb_o_ciphertext[448];
assign   tb_o_tag_ready[449]                  =   1'b0;
assign   tb_o_tag[449]                        =   tb_o_tag[448];

// CLK no. 450/1240
// *************************************************
assign   tb_i_valid[450]                      =   1'b0;
assign   tb_i_reset[450]                      =   1'b0;
assign   tb_i_sop[450]                        =   1'b0;
assign   tb_i_key_update[450]                 =   1'b0;
assign   tb_i_key[450]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[450]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[450]               =   1'b0;
assign   tb_i_rf_static_encrypt[450]          =   1'b1;
assign   tb_i_clear_fault_flags[450]          =   1'b0;
assign   tb_i_rf_static_aad_length[450]       =   64'h0000000000000100;
assign   tb_i_aad[450]                        =   tb_i_aad[449];
assign   tb_i_rf_static_plaintext_length[450] =   64'h0000000000000280;
assign   tb_i_plaintext[450]                  =   tb_i_plaintext[449];
assign   tb_o_valid[450]                      =   1'b0;
assign   tb_o_sop[450]                        =   1'b0;
assign   tb_o_ciphertext[450]                 =   tb_o_ciphertext[449];
assign   tb_o_tag_ready[450]                  =   1'b0;
assign   tb_o_tag[450]                        =   tb_o_tag[449];

// CLK no. 451/1240
// *************************************************
assign   tb_i_valid[451]                      =   1'b0;
assign   tb_i_reset[451]                      =   1'b0;
assign   tb_i_sop[451]                        =   1'b0;
assign   tb_i_key_update[451]                 =   1'b0;
assign   tb_i_key[451]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[451]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[451]               =   1'b0;
assign   tb_i_rf_static_encrypt[451]          =   1'b1;
assign   tb_i_clear_fault_flags[451]          =   1'b0;
assign   tb_i_rf_static_aad_length[451]       =   64'h0000000000000100;
assign   tb_i_aad[451]                        =   tb_i_aad[450];
assign   tb_i_rf_static_plaintext_length[451] =   64'h0000000000000280;
assign   tb_i_plaintext[451]                  =   tb_i_plaintext[450];
assign   tb_o_valid[451]                      =   1'b0;
assign   tb_o_sop[451]                        =   1'b0;
assign   tb_o_ciphertext[451]                 =   tb_o_ciphertext[450];
assign   tb_o_tag_ready[451]                  =   1'b0;
assign   tb_o_tag[451]                        =   tb_o_tag[450];

// CLK no. 452/1240
// *************************************************
assign   tb_i_valid[452]                      =   1'b0;
assign   tb_i_reset[452]                      =   1'b0;
assign   tb_i_sop[452]                        =   1'b0;
assign   tb_i_key_update[452]                 =   1'b0;
assign   tb_i_key[452]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[452]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[452]               =   1'b0;
assign   tb_i_rf_static_encrypt[452]          =   1'b1;
assign   tb_i_clear_fault_flags[452]          =   1'b0;
assign   tb_i_rf_static_aad_length[452]       =   64'h0000000000000100;
assign   tb_i_aad[452]                        =   tb_i_aad[451];
assign   tb_i_rf_static_plaintext_length[452] =   64'h0000000000000280;
assign   tb_i_plaintext[452]                  =   tb_i_plaintext[451];
assign   tb_o_valid[452]                      =   1'b0;
assign   tb_o_sop[452]                        =   1'b0;
assign   tb_o_ciphertext[452]                 =   tb_o_ciphertext[451];
assign   tb_o_tag_ready[452]                  =   1'b0;
assign   tb_o_tag[452]                        =   tb_o_tag[451];

// CLK no. 453/1240
// *************************************************
assign   tb_i_valid[453]                      =   1'b0;
assign   tb_i_reset[453]                      =   1'b0;
assign   tb_i_sop[453]                        =   1'b0;
assign   tb_i_key_update[453]                 =   1'b0;
assign   tb_i_key[453]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[453]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[453]               =   1'b0;
assign   tb_i_rf_static_encrypt[453]          =   1'b1;
assign   tb_i_clear_fault_flags[453]          =   1'b0;
assign   tb_i_rf_static_aad_length[453]       =   64'h0000000000000100;
assign   tb_i_aad[453]                        =   tb_i_aad[452];
assign   tb_i_rf_static_plaintext_length[453] =   64'h0000000000000280;
assign   tb_i_plaintext[453]                  =   tb_i_plaintext[452];
assign   tb_o_valid[453]                      =   1'b0;
assign   tb_o_sop[453]                        =   1'b0;
assign   tb_o_ciphertext[453]                 =   tb_o_ciphertext[452];
assign   tb_o_tag_ready[453]                  =   1'b0;
assign   tb_o_tag[453]                        =   tb_o_tag[452];

// CLK no. 454/1240
// *************************************************
assign   tb_i_valid[454]                      =   1'b0;
assign   tb_i_reset[454]                      =   1'b0;
assign   tb_i_sop[454]                        =   1'b0;
assign   tb_i_key_update[454]                 =   1'b0;
assign   tb_i_key[454]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[454]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[454]               =   1'b0;
assign   tb_i_rf_static_encrypt[454]          =   1'b1;
assign   tb_i_clear_fault_flags[454]          =   1'b0;
assign   tb_i_rf_static_aad_length[454]       =   64'h0000000000000100;
assign   tb_i_aad[454]                        =   tb_i_aad[453];
assign   tb_i_rf_static_plaintext_length[454] =   64'h0000000000000280;
assign   tb_i_plaintext[454]                  =   tb_i_plaintext[453];
assign   tb_o_valid[454]                      =   1'b0;
assign   tb_o_sop[454]                        =   1'b0;
assign   tb_o_ciphertext[454]                 =   tb_o_ciphertext[453];
assign   tb_o_tag_ready[454]                  =   1'b0;
assign   tb_o_tag[454]                        =   tb_o_tag[453];

// CLK no. 455/1240
// *************************************************
assign   tb_i_valid[455]                      =   1'b0;
assign   tb_i_reset[455]                      =   1'b0;
assign   tb_i_sop[455]                        =   1'b0;
assign   tb_i_key_update[455]                 =   1'b0;
assign   tb_i_key[455]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[455]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[455]               =   1'b0;
assign   tb_i_rf_static_encrypt[455]          =   1'b1;
assign   tb_i_clear_fault_flags[455]          =   1'b0;
assign   tb_i_rf_static_aad_length[455]       =   64'h0000000000000100;
assign   tb_i_aad[455]                        =   tb_i_aad[454];
assign   tb_i_rf_static_plaintext_length[455] =   64'h0000000000000280;
assign   tb_i_plaintext[455]                  =   tb_i_plaintext[454];
assign   tb_o_valid[455]                      =   1'b0;
assign   tb_o_sop[455]                        =   1'b0;
assign   tb_o_ciphertext[455]                 =   tb_o_ciphertext[454];
assign   tb_o_tag_ready[455]                  =   1'b0;
assign   tb_o_tag[455]                        =   tb_o_tag[454];

// CLK no. 456/1240
// *************************************************
assign   tb_i_valid[456]                      =   1'b0;
assign   tb_i_reset[456]                      =   1'b0;
assign   tb_i_sop[456]                        =   1'b0;
assign   tb_i_key_update[456]                 =   1'b0;
assign   tb_i_key[456]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[456]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[456]               =   1'b0;
assign   tb_i_rf_static_encrypt[456]          =   1'b1;
assign   tb_i_clear_fault_flags[456]          =   1'b0;
assign   tb_i_rf_static_aad_length[456]       =   64'h0000000000000100;
assign   tb_i_aad[456]                        =   tb_i_aad[455];
assign   tb_i_rf_static_plaintext_length[456] =   64'h0000000000000280;
assign   tb_i_plaintext[456]                  =   tb_i_plaintext[455];
assign   tb_o_valid[456]                      =   1'b0;
assign   tb_o_sop[456]                        =   1'b0;
assign   tb_o_ciphertext[456]                 =   tb_o_ciphertext[455];
assign   tb_o_tag_ready[456]                  =   1'b0;
assign   tb_o_tag[456]                        =   tb_o_tag[455];

// CLK no. 457/1240
// *************************************************
assign   tb_i_valid[457]                      =   1'b0;
assign   tb_i_reset[457]                      =   1'b0;
assign   tb_i_sop[457]                        =   1'b0;
assign   tb_i_key_update[457]                 =   1'b0;
assign   tb_i_key[457]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[457]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[457]               =   1'b0;
assign   tb_i_rf_static_encrypt[457]          =   1'b1;
assign   tb_i_clear_fault_flags[457]          =   1'b0;
assign   tb_i_rf_static_aad_length[457]       =   64'h0000000000000100;
assign   tb_i_aad[457]                        =   tb_i_aad[456];
assign   tb_i_rf_static_plaintext_length[457] =   64'h0000000000000280;
assign   tb_i_plaintext[457]                  =   tb_i_plaintext[456];
assign   tb_o_valid[457]                      =   1'b0;
assign   tb_o_sop[457]                        =   1'b0;
assign   tb_o_ciphertext[457]                 =   tb_o_ciphertext[456];
assign   tb_o_tag_ready[457]                  =   1'b0;
assign   tb_o_tag[457]                        =   tb_o_tag[456];

// CLK no. 458/1240
// *************************************************
assign   tb_i_valid[458]                      =   1'b0;
assign   tb_i_reset[458]                      =   1'b0;
assign   tb_i_sop[458]                        =   1'b0;
assign   tb_i_key_update[458]                 =   1'b0;
assign   tb_i_key[458]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[458]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[458]               =   1'b0;
assign   tb_i_rf_static_encrypt[458]          =   1'b1;
assign   tb_i_clear_fault_flags[458]          =   1'b0;
assign   tb_i_rf_static_aad_length[458]       =   64'h0000000000000100;
assign   tb_i_aad[458]                        =   tb_i_aad[457];
assign   tb_i_rf_static_plaintext_length[458] =   64'h0000000000000280;
assign   tb_i_plaintext[458]                  =   tb_i_plaintext[457];
assign   tb_o_valid[458]                      =   1'b0;
assign   tb_o_sop[458]                        =   1'b0;
assign   tb_o_ciphertext[458]                 =   tb_o_ciphertext[457];
assign   tb_o_tag_ready[458]                  =   1'b0;
assign   tb_o_tag[458]                        =   tb_o_tag[457];

// CLK no. 459/1240
// *************************************************
assign   tb_i_valid[459]                      =   1'b0;
assign   tb_i_reset[459]                      =   1'b0;
assign   tb_i_sop[459]                        =   1'b0;
assign   tb_i_key_update[459]                 =   1'b0;
assign   tb_i_key[459]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[459]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[459]               =   1'b0;
assign   tb_i_rf_static_encrypt[459]          =   1'b1;
assign   tb_i_clear_fault_flags[459]          =   1'b0;
assign   tb_i_rf_static_aad_length[459]       =   64'h0000000000000100;
assign   tb_i_aad[459]                        =   tb_i_aad[458];
assign   tb_i_rf_static_plaintext_length[459] =   64'h0000000000000280;
assign   tb_i_plaintext[459]                  =   tb_i_plaintext[458];
assign   tb_o_valid[459]                      =   1'b0;
assign   tb_o_sop[459]                        =   1'b0;
assign   tb_o_ciphertext[459]                 =   tb_o_ciphertext[458];
assign   tb_o_tag_ready[459]                  =   1'b0;
assign   tb_o_tag[459]                        =   tb_o_tag[458];

// CLK no. 460/1240
// *************************************************
assign   tb_i_valid[460]                      =   1'b0;
assign   tb_i_reset[460]                      =   1'b0;
assign   tb_i_sop[460]                        =   1'b0;
assign   tb_i_key_update[460]                 =   1'b0;
assign   tb_i_key[460]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[460]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[460]               =   1'b0;
assign   tb_i_rf_static_encrypt[460]          =   1'b1;
assign   tb_i_clear_fault_flags[460]          =   1'b0;
assign   tb_i_rf_static_aad_length[460]       =   64'h0000000000000100;
assign   tb_i_aad[460]                        =   tb_i_aad[459];
assign   tb_i_rf_static_plaintext_length[460] =   64'h0000000000000280;
assign   tb_i_plaintext[460]                  =   tb_i_plaintext[459];
assign   tb_o_valid[460]                      =   1'b1;
assign   tb_o_sop[460]                        =   1'b1;
assign   tb_o_ciphertext[460]                 =   256'ha714bfe727684d33021a0e7aa2b1e0f1510aa248591f6022d1e162c4eef39d70;
assign   tb_o_tag_ready[460]                  =   1'b0;
assign   tb_o_tag[460]                        =   tb_o_tag[459];

// CLK no. 461/1240
// *************************************************
assign   tb_i_valid[461]                      =   1'b0;
assign   tb_i_reset[461]                      =   1'b0;
assign   tb_i_sop[461]                        =   1'b0;
assign   tb_i_key_update[461]                 =   1'b0;
assign   tb_i_key[461]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[461]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[461]               =   1'b0;
assign   tb_i_rf_static_encrypt[461]          =   1'b1;
assign   tb_i_clear_fault_flags[461]          =   1'b0;
assign   tb_i_rf_static_aad_length[461]       =   64'h0000000000000100;
assign   tb_i_aad[461]                        =   tb_i_aad[460];
assign   tb_i_rf_static_plaintext_length[461] =   64'h0000000000000280;
assign   tb_i_plaintext[461]                  =   tb_i_plaintext[460];
assign   tb_o_valid[461]                      =   1'b1;
assign   tb_o_sop[461]                        =   1'b0;
assign   tb_o_ciphertext[461]                 =   256'ha36a04853da40adafc84080de632c73169ed9c52f41da327de31416269796d96;
assign   tb_o_tag_ready[461]                  =   1'b0;
assign   tb_o_tag[461]                        =   tb_o_tag[460];

// CLK no. 462/1240
// *************************************************
assign   tb_i_valid[462]                      =   1'b0;
assign   tb_i_reset[462]                      =   1'b0;
assign   tb_i_sop[462]                        =   1'b0;
assign   tb_i_key_update[462]                 =   1'b0;
assign   tb_i_key[462]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[462]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[462]               =   1'b0;
assign   tb_i_rf_static_encrypt[462]          =   1'b1;
assign   tb_i_clear_fault_flags[462]          =   1'b0;
assign   tb_i_rf_static_aad_length[462]       =   64'h0000000000000100;
assign   tb_i_aad[462]                        =   tb_i_aad[461];
assign   tb_i_rf_static_plaintext_length[462] =   64'h0000000000000280;
assign   tb_i_plaintext[462]                  =   tb_i_plaintext[461];
assign   tb_o_valid[462]                      =   1'b1;
assign   tb_o_sop[462]                        =   1'b0;
assign   tb_o_ciphertext[462]                 =   256'ha5f7ea767dbad0fce2723e314cd5eb64;
assign   tb_o_tag_ready[462]                  =   1'b0;
assign   tb_o_tag[462]                        =   tb_o_tag[461];

// CLK no. 463/1240
// *************************************************
assign   tb_i_valid[463]                      =   1'b0;
assign   tb_i_reset[463]                      =   1'b0;
assign   tb_i_sop[463]                        =   1'b0;
assign   tb_i_key_update[463]                 =   1'b0;
assign   tb_i_key[463]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[463]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[463]               =   1'b0;
assign   tb_i_rf_static_encrypt[463]          =   1'b1;
assign   tb_i_clear_fault_flags[463]          =   1'b0;
assign   tb_i_rf_static_aad_length[463]       =   64'h0000000000000100;
assign   tb_i_aad[463]                        =   tb_i_aad[462];
assign   tb_i_rf_static_plaintext_length[463] =   64'h0000000000000280;
assign   tb_i_plaintext[463]                  =   tb_i_plaintext[462];
assign   tb_o_valid[463]                      =   1'b0;
assign   tb_o_sop[463]                        =   1'b0;
assign   tb_o_ciphertext[463]                 =   tb_o_ciphertext[462];
assign   tb_o_tag_ready[463]                  =   1'b0;
assign   tb_o_tag[463]                        =   tb_o_tag[462];

// CLK no. 464/1240
// *************************************************
assign   tb_i_valid[464]                      =   1'b0;
assign   tb_i_reset[464]                      =   1'b0;
assign   tb_i_sop[464]                        =   1'b0;
assign   tb_i_key_update[464]                 =   1'b0;
assign   tb_i_key[464]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[464]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[464]               =   1'b0;
assign   tb_i_rf_static_encrypt[464]          =   1'b1;
assign   tb_i_clear_fault_flags[464]          =   1'b0;
assign   tb_i_rf_static_aad_length[464]       =   64'h0000000000000100;
assign   tb_i_aad[464]                        =   tb_i_aad[463];
assign   tb_i_rf_static_plaintext_length[464] =   64'h0000000000000280;
assign   tb_i_plaintext[464]                  =   tb_i_plaintext[463];
assign   tb_o_valid[464]                      =   1'b0;
assign   tb_o_sop[464]                        =   1'b0;
assign   tb_o_ciphertext[464]                 =   tb_o_ciphertext[463];
assign   tb_o_tag_ready[464]                  =   1'b0;
assign   tb_o_tag[464]                        =   tb_o_tag[463];

// CLK no. 465/1240
// *************************************************
assign   tb_i_valid[465]                      =   1'b0;
assign   tb_i_reset[465]                      =   1'b0;
assign   tb_i_sop[465]                        =   1'b0;
assign   tb_i_key_update[465]                 =   1'b0;
assign   tb_i_key[465]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[465]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[465]               =   1'b0;
assign   tb_i_rf_static_encrypt[465]          =   1'b1;
assign   tb_i_clear_fault_flags[465]          =   1'b0;
assign   tb_i_rf_static_aad_length[465]       =   64'h0000000000000100;
assign   tb_i_aad[465]                        =   tb_i_aad[464];
assign   tb_i_rf_static_plaintext_length[465] =   64'h0000000000000280;
assign   tb_i_plaintext[465]                  =   tb_i_plaintext[464];
assign   tb_o_valid[465]                      =   1'b0;
assign   tb_o_sop[465]                        =   1'b0;
assign   tb_o_ciphertext[465]                 =   tb_o_ciphertext[464];
assign   tb_o_tag_ready[465]                  =   1'b0;
assign   tb_o_tag[465]                        =   tb_o_tag[464];

// CLK no. 466/1240
// *************************************************
assign   tb_i_valid[466]                      =   1'b0;
assign   tb_i_reset[466]                      =   1'b0;
assign   tb_i_sop[466]                        =   1'b0;
assign   tb_i_key_update[466]                 =   1'b0;
assign   tb_i_key[466]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[466]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[466]               =   1'b0;
assign   tb_i_rf_static_encrypt[466]          =   1'b1;
assign   tb_i_clear_fault_flags[466]          =   1'b0;
assign   tb_i_rf_static_aad_length[466]       =   64'h0000000000000100;
assign   tb_i_aad[466]                        =   tb_i_aad[465];
assign   tb_i_rf_static_plaintext_length[466] =   64'h0000000000000280;
assign   tb_i_plaintext[466]                  =   tb_i_plaintext[465];
assign   tb_o_valid[466]                      =   1'b0;
assign   tb_o_sop[466]                        =   1'b0;
assign   tb_o_ciphertext[466]                 =   tb_o_ciphertext[465];
assign   tb_o_tag_ready[466]                  =   1'b0;
assign   tb_o_tag[466]                        =   tb_o_tag[465];

// CLK no. 467/1240
// *************************************************
assign   tb_i_valid[467]                      =   1'b0;
assign   tb_i_reset[467]                      =   1'b0;
assign   tb_i_sop[467]                        =   1'b0;
assign   tb_i_key_update[467]                 =   1'b0;
assign   tb_i_key[467]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[467]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[467]               =   1'b0;
assign   tb_i_rf_static_encrypt[467]          =   1'b1;
assign   tb_i_clear_fault_flags[467]          =   1'b0;
assign   tb_i_rf_static_aad_length[467]       =   64'h0000000000000100;
assign   tb_i_aad[467]                        =   tb_i_aad[466];
assign   tb_i_rf_static_plaintext_length[467] =   64'h0000000000000280;
assign   tb_i_plaintext[467]                  =   tb_i_plaintext[466];
assign   tb_o_valid[467]                      =   1'b0;
assign   tb_o_sop[467]                        =   1'b0;
assign   tb_o_ciphertext[467]                 =   tb_o_ciphertext[466];
assign   tb_o_tag_ready[467]                  =   1'b0;
assign   tb_o_tag[467]                        =   tb_o_tag[466];

// CLK no. 468/1240
// *************************************************
assign   tb_i_valid[468]                      =   1'b0;
assign   tb_i_reset[468]                      =   1'b0;
assign   tb_i_sop[468]                        =   1'b0;
assign   tb_i_key_update[468]                 =   1'b0;
assign   tb_i_key[468]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[468]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[468]               =   1'b0;
assign   tb_i_rf_static_encrypt[468]          =   1'b1;
assign   tb_i_clear_fault_flags[468]          =   1'b0;
assign   tb_i_rf_static_aad_length[468]       =   64'h0000000000000100;
assign   tb_i_aad[468]                        =   tb_i_aad[467];
assign   tb_i_rf_static_plaintext_length[468] =   64'h0000000000000280;
assign   tb_i_plaintext[468]                  =   tb_i_plaintext[467];
assign   tb_o_valid[468]                      =   1'b0;
assign   tb_o_sop[468]                        =   1'b0;
assign   tb_o_ciphertext[468]                 =   tb_o_ciphertext[467];
assign   tb_o_tag_ready[468]                  =   1'b0;
assign   tb_o_tag[468]                        =   tb_o_tag[467];

// CLK no. 469/1240
// *************************************************
assign   tb_i_valid[469]                      =   1'b0;
assign   tb_i_reset[469]                      =   1'b0;
assign   tb_i_sop[469]                        =   1'b0;
assign   tb_i_key_update[469]                 =   1'b0;
assign   tb_i_key[469]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[469]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[469]               =   1'b0;
assign   tb_i_rf_static_encrypt[469]          =   1'b1;
assign   tb_i_clear_fault_flags[469]          =   1'b0;
assign   tb_i_rf_static_aad_length[469]       =   64'h0000000000000100;
assign   tb_i_aad[469]                        =   tb_i_aad[468];
assign   tb_i_rf_static_plaintext_length[469] =   64'h0000000000000280;
assign   tb_i_plaintext[469]                  =   tb_i_plaintext[468];
assign   tb_o_valid[469]                      =   1'b0;
assign   tb_o_sop[469]                        =   1'b0;
assign   tb_o_ciphertext[469]                 =   tb_o_ciphertext[468];
assign   tb_o_tag_ready[469]                  =   1'b0;
assign   tb_o_tag[469]                        =   tb_o_tag[468];

// CLK no. 470/1240
// *************************************************
assign   tb_i_valid[470]                      =   1'b0;
assign   tb_i_reset[470]                      =   1'b0;
assign   tb_i_sop[470]                        =   1'b0;
assign   tb_i_key_update[470]                 =   1'b0;
assign   tb_i_key[470]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[470]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[470]               =   1'b0;
assign   tb_i_rf_static_encrypt[470]          =   1'b1;
assign   tb_i_clear_fault_flags[470]          =   1'b0;
assign   tb_i_rf_static_aad_length[470]       =   64'h0000000000000100;
assign   tb_i_aad[470]                        =   tb_i_aad[469];
assign   tb_i_rf_static_plaintext_length[470] =   64'h0000000000000280;
assign   tb_i_plaintext[470]                  =   tb_i_plaintext[469];
assign   tb_o_valid[470]                      =   1'b0;
assign   tb_o_sop[470]                        =   1'b0;
assign   tb_o_ciphertext[470]                 =   tb_o_ciphertext[469];
assign   tb_o_tag_ready[470]                  =   1'b1;
assign   tb_o_tag[470]                        =   128'h5b0e3365a64e77debd90ff20e3729bfe;

// CLK no. 471/1240
// *************************************************
assign   tb_i_valid[471]                      =   1'b0;
assign   tb_i_reset[471]                      =   1'b0;
assign   tb_i_sop[471]                        =   1'b0;
assign   tb_i_key_update[471]                 =   1'b0;
assign   tb_i_key[471]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[471]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[471]               =   1'b0;
assign   tb_i_rf_static_encrypt[471]          =   1'b1;
assign   tb_i_clear_fault_flags[471]          =   1'b0;
assign   tb_i_rf_static_aad_length[471]       =   64'h0000000000000100;
assign   tb_i_aad[471]                        =   tb_i_aad[470];
assign   tb_i_rf_static_plaintext_length[471] =   64'h0000000000000280;
assign   tb_i_plaintext[471]                  =   tb_i_plaintext[470];
assign   tb_o_valid[471]                      =   1'b0;
assign   tb_o_sop[471]                        =   1'b0;
assign   tb_o_ciphertext[471]                 =   tb_o_ciphertext[470];
assign   tb_o_tag_ready[471]                  =   1'b0;
assign   tb_o_tag[471]                        =   tb_o_tag[470];

// CLK no. 472/1240
// *************************************************
assign   tb_i_valid[472]                      =   1'b0;
assign   tb_i_reset[472]                      =   1'b0;
assign   tb_i_sop[472]                        =   1'b0;
assign   tb_i_key_update[472]                 =   1'b0;
assign   tb_i_key[472]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[472]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[472]               =   1'b0;
assign   tb_i_rf_static_encrypt[472]          =   1'b1;
assign   tb_i_clear_fault_flags[472]          =   1'b0;
assign   tb_i_rf_static_aad_length[472]       =   64'h0000000000000100;
assign   tb_i_aad[472]                        =   tb_i_aad[471];
assign   tb_i_rf_static_plaintext_length[472] =   64'h0000000000000280;
assign   tb_i_plaintext[472]                  =   tb_i_plaintext[471];
assign   tb_o_valid[472]                      =   1'b0;
assign   tb_o_sop[472]                        =   1'b0;
assign   tb_o_ciphertext[472]                 =   tb_o_ciphertext[471];
assign   tb_o_tag_ready[472]                  =   1'b0;
assign   tb_o_tag[472]                        =   tb_o_tag[471];

// CLK no. 473/1240
// *************************************************
assign   tb_i_valid[473]                      =   1'b0;
assign   tb_i_reset[473]                      =   1'b0;
assign   tb_i_sop[473]                        =   1'b1;
assign   tb_i_key_update[473]                 =   1'b0;
assign   tb_i_key[473]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[473]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[473]               =   1'b0;
assign   tb_i_rf_static_encrypt[473]          =   1'b1;
assign   tb_i_clear_fault_flags[473]          =   1'b0;
assign   tb_i_rf_static_aad_length[473]       =   64'h0000000000000100;
assign   tb_i_aad[473]                        =   tb_i_aad[472];
assign   tb_i_rf_static_plaintext_length[473] =   64'h0000000000000280;
assign   tb_i_plaintext[473]                  =   tb_i_plaintext[472];
assign   tb_o_valid[473]                      =   1'b0;
assign   tb_o_sop[473]                        =   1'b0;
assign   tb_o_ciphertext[473]                 =   tb_o_ciphertext[472];
assign   tb_o_tag_ready[473]                  =   1'b0;
assign   tb_o_tag[473]                        =   tb_o_tag[472];

// CLK no. 474/1240
// *************************************************
assign   tb_i_valid[474]                      =   1'b1;
assign   tb_i_reset[474]                      =   1'b0;
assign   tb_i_sop[474]                        =   1'b0;
assign   tb_i_key_update[474]                 =   1'b0;
assign   tb_i_key[474]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[474]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[474]               =   1'b0;
assign   tb_i_rf_static_encrypt[474]          =   1'b1;
assign   tb_i_clear_fault_flags[474]          =   1'b0;
assign   tb_i_rf_static_aad_length[474]       =   64'h0000000000000100;
assign   tb_i_aad[474]                        =   256'h50abe8ec8bd84ad3e87e22150fef13b168aadb6e2dc3feb58a03f4d92b1a161e;
assign   tb_i_rf_static_plaintext_length[474] =   64'h0000000000000280;
assign   tb_i_plaintext[474]                  =   tb_i_plaintext[473];
assign   tb_o_valid[474]                      =   1'b0;
assign   tb_o_sop[474]                        =   1'b0;
assign   tb_o_ciphertext[474]                 =   tb_o_ciphertext[473];
assign   tb_o_tag_ready[474]                  =   1'b0;
assign   tb_o_tag[474]                        =   tb_o_tag[473];

// CLK no. 475/1240
// *************************************************
assign   tb_i_valid[475]                      =   1'b1;
assign   tb_i_reset[475]                      =   1'b0;
assign   tb_i_sop[475]                        =   1'b0;
assign   tb_i_key_update[475]                 =   1'b0;
assign   tb_i_key[475]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[475]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[475]               =   1'b0;
assign   tb_i_rf_static_encrypt[475]          =   1'b1;
assign   tb_i_clear_fault_flags[475]          =   1'b0;
assign   tb_i_rf_static_aad_length[475]       =   64'h0000000000000100;
assign   tb_i_aad[475]                        =   tb_i_aad[474];
assign   tb_i_rf_static_plaintext_length[475] =   64'h0000000000000280;
assign   tb_i_plaintext[475]                  =   256'h9af988663fae50f8c15c7026c7aecc2d3a7e850ab68893f84fb087490c18b338;
assign   tb_o_valid[475]                      =   1'b0;
assign   tb_o_sop[475]                        =   1'b0;
assign   tb_o_ciphertext[475]                 =   tb_o_ciphertext[474];
assign   tb_o_tag_ready[475]                  =   1'b0;
assign   tb_o_tag[475]                        =   tb_o_tag[474];

// CLK no. 476/1240
// *************************************************
assign   tb_i_valid[476]                      =   1'b1;
assign   tb_i_reset[476]                      =   1'b0;
assign   tb_i_sop[476]                        =   1'b0;
assign   tb_i_key_update[476]                 =   1'b0;
assign   tb_i_key[476]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[476]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[476]               =   1'b0;
assign   tb_i_rf_static_encrypt[476]          =   1'b1;
assign   tb_i_clear_fault_flags[476]          =   1'b0;
assign   tb_i_rf_static_aad_length[476]       =   64'h0000000000000100;
assign   tb_i_aad[476]                        =   tb_i_aad[475];
assign   tb_i_rf_static_plaintext_length[476] =   64'h0000000000000280;
assign   tb_i_plaintext[476]                  =   256'h0a2ddcf2148b86e1a9396fee6d5568f799161cf8c45f2eea171a34d281493496;
assign   tb_o_valid[476]                      =   1'b0;
assign   tb_o_sop[476]                        =   1'b0;
assign   tb_o_ciphertext[476]                 =   tb_o_ciphertext[475];
assign   tb_o_tag_ready[476]                  =   1'b0;
assign   tb_o_tag[476]                        =   tb_o_tag[475];

// CLK no. 477/1240
// *************************************************
assign   tb_i_valid[477]                      =   1'b1;
assign   tb_i_reset[477]                      =   1'b0;
assign   tb_i_sop[477]                        =   1'b0;
assign   tb_i_key_update[477]                 =   1'b0;
assign   tb_i_key[477]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[477]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[477]               =   1'b0;
assign   tb_i_rf_static_encrypt[477]          =   1'b1;
assign   tb_i_clear_fault_flags[477]          =   1'b0;
assign   tb_i_rf_static_aad_length[477]       =   64'h0000000000000100;
assign   tb_i_aad[477]                        =   tb_i_aad[476];
assign   tb_i_rf_static_plaintext_length[477] =   64'h0000000000000280;
assign   tb_i_plaintext[477]                  =   256'ha6ae802d649ff8a1350837c2090bd74a;
assign   tb_o_valid[477]                      =   1'b0;
assign   tb_o_sop[477]                        =   1'b0;
assign   tb_o_ciphertext[477]                 =   tb_o_ciphertext[476];
assign   tb_o_tag_ready[477]                  =   1'b0;
assign   tb_o_tag[477]                        =   tb_o_tag[476];

// CLK no. 478/1240
// *************************************************
assign   tb_i_valid[478]                      =   1'b0;
assign   tb_i_reset[478]                      =   1'b0;
assign   tb_i_sop[478]                        =   1'b0;
assign   tb_i_key_update[478]                 =   1'b0;
assign   tb_i_key[478]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[478]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[478]               =   1'b0;
assign   tb_i_rf_static_encrypt[478]          =   1'b1;
assign   tb_i_clear_fault_flags[478]          =   1'b0;
assign   tb_i_rf_static_aad_length[478]       =   64'h0000000000000100;
assign   tb_i_aad[478]                        =   tb_i_aad[477];
assign   tb_i_rf_static_plaintext_length[478] =   64'h0000000000000280;
assign   tb_i_plaintext[478]                  =   tb_i_plaintext[477];
assign   tb_o_valid[478]                      =   1'b0;
assign   tb_o_sop[478]                        =   1'b0;
assign   tb_o_ciphertext[478]                 =   tb_o_ciphertext[477];
assign   tb_o_tag_ready[478]                  =   1'b0;
assign   tb_o_tag[478]                        =   tb_o_tag[477];

// CLK no. 479/1240
// *************************************************
assign   tb_i_valid[479]                      =   1'b0;
assign   tb_i_reset[479]                      =   1'b0;
assign   tb_i_sop[479]                        =   1'b0;
assign   tb_i_key_update[479]                 =   1'b0;
assign   tb_i_key[479]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[479]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[479]               =   1'b0;
assign   tb_i_rf_static_encrypt[479]          =   1'b1;
assign   tb_i_clear_fault_flags[479]          =   1'b0;
assign   tb_i_rf_static_aad_length[479]       =   64'h0000000000000100;
assign   tb_i_aad[479]                        =   tb_i_aad[478];
assign   tb_i_rf_static_plaintext_length[479] =   64'h0000000000000280;
assign   tb_i_plaintext[479]                  =   tb_i_plaintext[478];
assign   tb_o_valid[479]                      =   1'b0;
assign   tb_o_sop[479]                        =   1'b0;
assign   tb_o_ciphertext[479]                 =   tb_o_ciphertext[478];
assign   tb_o_tag_ready[479]                  =   1'b0;
assign   tb_o_tag[479]                        =   tb_o_tag[478];

// CLK no. 480/1240
// *************************************************
assign   tb_i_valid[480]                      =   1'b0;
assign   tb_i_reset[480]                      =   1'b0;
assign   tb_i_sop[480]                        =   1'b0;
assign   tb_i_key_update[480]                 =   1'b0;
assign   tb_i_key[480]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[480]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[480]               =   1'b0;
assign   tb_i_rf_static_encrypt[480]          =   1'b1;
assign   tb_i_clear_fault_flags[480]          =   1'b0;
assign   tb_i_rf_static_aad_length[480]       =   64'h0000000000000100;
assign   tb_i_aad[480]                        =   tb_i_aad[479];
assign   tb_i_rf_static_plaintext_length[480] =   64'h0000000000000280;
assign   tb_i_plaintext[480]                  =   tb_i_plaintext[479];
assign   tb_o_valid[480]                      =   1'b0;
assign   tb_o_sop[480]                        =   1'b0;
assign   tb_o_ciphertext[480]                 =   tb_o_ciphertext[479];
assign   tb_o_tag_ready[480]                  =   1'b0;
assign   tb_o_tag[480]                        =   tb_o_tag[479];

// CLK no. 481/1240
// *************************************************
assign   tb_i_valid[481]                      =   1'b0;
assign   tb_i_reset[481]                      =   1'b0;
assign   tb_i_sop[481]                        =   1'b0;
assign   tb_i_key_update[481]                 =   1'b0;
assign   tb_i_key[481]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[481]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[481]               =   1'b0;
assign   tb_i_rf_static_encrypt[481]          =   1'b1;
assign   tb_i_clear_fault_flags[481]          =   1'b0;
assign   tb_i_rf_static_aad_length[481]       =   64'h0000000000000100;
assign   tb_i_aad[481]                        =   tb_i_aad[480];
assign   tb_i_rf_static_plaintext_length[481] =   64'h0000000000000280;
assign   tb_i_plaintext[481]                  =   tb_i_plaintext[480];
assign   tb_o_valid[481]                      =   1'b0;
assign   tb_o_sop[481]                        =   1'b0;
assign   tb_o_ciphertext[481]                 =   tb_o_ciphertext[480];
assign   tb_o_tag_ready[481]                  =   1'b0;
assign   tb_o_tag[481]                        =   tb_o_tag[480];

// CLK no. 482/1240
// *************************************************
assign   tb_i_valid[482]                      =   1'b0;
assign   tb_i_reset[482]                      =   1'b0;
assign   tb_i_sop[482]                        =   1'b0;
assign   tb_i_key_update[482]                 =   1'b0;
assign   tb_i_key[482]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[482]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[482]               =   1'b0;
assign   tb_i_rf_static_encrypt[482]          =   1'b1;
assign   tb_i_clear_fault_flags[482]          =   1'b0;
assign   tb_i_rf_static_aad_length[482]       =   64'h0000000000000100;
assign   tb_i_aad[482]                        =   tb_i_aad[481];
assign   tb_i_rf_static_plaintext_length[482] =   64'h0000000000000280;
assign   tb_i_plaintext[482]                  =   tb_i_plaintext[481];
assign   tb_o_valid[482]                      =   1'b0;
assign   tb_o_sop[482]                        =   1'b0;
assign   tb_o_ciphertext[482]                 =   tb_o_ciphertext[481];
assign   tb_o_tag_ready[482]                  =   1'b0;
assign   tb_o_tag[482]                        =   tb_o_tag[481];

// CLK no. 483/1240
// *************************************************
assign   tb_i_valid[483]                      =   1'b0;
assign   tb_i_reset[483]                      =   1'b0;
assign   tb_i_sop[483]                        =   1'b0;
assign   tb_i_key_update[483]                 =   1'b0;
assign   tb_i_key[483]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[483]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[483]               =   1'b0;
assign   tb_i_rf_static_encrypt[483]          =   1'b1;
assign   tb_i_clear_fault_flags[483]          =   1'b0;
assign   tb_i_rf_static_aad_length[483]       =   64'h0000000000000100;
assign   tb_i_aad[483]                        =   tb_i_aad[482];
assign   tb_i_rf_static_plaintext_length[483] =   64'h0000000000000280;
assign   tb_i_plaintext[483]                  =   tb_i_plaintext[482];
assign   tb_o_valid[483]                      =   1'b0;
assign   tb_o_sop[483]                        =   1'b0;
assign   tb_o_ciphertext[483]                 =   tb_o_ciphertext[482];
assign   tb_o_tag_ready[483]                  =   1'b0;
assign   tb_o_tag[483]                        =   tb_o_tag[482];

// CLK no. 484/1240
// *************************************************
assign   tb_i_valid[484]                      =   1'b0;
assign   tb_i_reset[484]                      =   1'b0;
assign   tb_i_sop[484]                        =   1'b0;
assign   tb_i_key_update[484]                 =   1'b0;
assign   tb_i_key[484]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[484]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[484]               =   1'b0;
assign   tb_i_rf_static_encrypt[484]          =   1'b1;
assign   tb_i_clear_fault_flags[484]          =   1'b0;
assign   tb_i_rf_static_aad_length[484]       =   64'h0000000000000100;
assign   tb_i_aad[484]                        =   tb_i_aad[483];
assign   tb_i_rf_static_plaintext_length[484] =   64'h0000000000000280;
assign   tb_i_plaintext[484]                  =   tb_i_plaintext[483];
assign   tb_o_valid[484]                      =   1'b0;
assign   tb_o_sop[484]                        =   1'b0;
assign   tb_o_ciphertext[484]                 =   tb_o_ciphertext[483];
assign   tb_o_tag_ready[484]                  =   1'b0;
assign   tb_o_tag[484]                        =   tb_o_tag[483];

// CLK no. 485/1240
// *************************************************
assign   tb_i_valid[485]                      =   1'b0;
assign   tb_i_reset[485]                      =   1'b0;
assign   tb_i_sop[485]                        =   1'b0;
assign   tb_i_key_update[485]                 =   1'b0;
assign   tb_i_key[485]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[485]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[485]               =   1'b0;
assign   tb_i_rf_static_encrypt[485]          =   1'b1;
assign   tb_i_clear_fault_flags[485]          =   1'b0;
assign   tb_i_rf_static_aad_length[485]       =   64'h0000000000000100;
assign   tb_i_aad[485]                        =   tb_i_aad[484];
assign   tb_i_rf_static_plaintext_length[485] =   64'h0000000000000280;
assign   tb_i_plaintext[485]                  =   tb_i_plaintext[484];
assign   tb_o_valid[485]                      =   1'b0;
assign   tb_o_sop[485]                        =   1'b0;
assign   tb_o_ciphertext[485]                 =   tb_o_ciphertext[484];
assign   tb_o_tag_ready[485]                  =   1'b0;
assign   tb_o_tag[485]                        =   tb_o_tag[484];

// CLK no. 486/1240
// *************************************************
assign   tb_i_valid[486]                      =   1'b0;
assign   tb_i_reset[486]                      =   1'b0;
assign   tb_i_sop[486]                        =   1'b0;
assign   tb_i_key_update[486]                 =   1'b0;
assign   tb_i_key[486]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[486]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[486]               =   1'b0;
assign   tb_i_rf_static_encrypt[486]          =   1'b1;
assign   tb_i_clear_fault_flags[486]          =   1'b0;
assign   tb_i_rf_static_aad_length[486]       =   64'h0000000000000100;
assign   tb_i_aad[486]                        =   tb_i_aad[485];
assign   tb_i_rf_static_plaintext_length[486] =   64'h0000000000000280;
assign   tb_i_plaintext[486]                  =   tb_i_plaintext[485];
assign   tb_o_valid[486]                      =   1'b0;
assign   tb_o_sop[486]                        =   1'b0;
assign   tb_o_ciphertext[486]                 =   tb_o_ciphertext[485];
assign   tb_o_tag_ready[486]                  =   1'b0;
assign   tb_o_tag[486]                        =   tb_o_tag[485];

// CLK no. 487/1240
// *************************************************
assign   tb_i_valid[487]                      =   1'b0;
assign   tb_i_reset[487]                      =   1'b0;
assign   tb_i_sop[487]                        =   1'b0;
assign   tb_i_key_update[487]                 =   1'b0;
assign   tb_i_key[487]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[487]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[487]               =   1'b0;
assign   tb_i_rf_static_encrypt[487]          =   1'b1;
assign   tb_i_clear_fault_flags[487]          =   1'b0;
assign   tb_i_rf_static_aad_length[487]       =   64'h0000000000000100;
assign   tb_i_aad[487]                        =   tb_i_aad[486];
assign   tb_i_rf_static_plaintext_length[487] =   64'h0000000000000280;
assign   tb_i_plaintext[487]                  =   tb_i_plaintext[486];
assign   tb_o_valid[487]                      =   1'b0;
assign   tb_o_sop[487]                        =   1'b0;
assign   tb_o_ciphertext[487]                 =   tb_o_ciphertext[486];
assign   tb_o_tag_ready[487]                  =   1'b0;
assign   tb_o_tag[487]                        =   tb_o_tag[486];

// CLK no. 488/1240
// *************************************************
assign   tb_i_valid[488]                      =   1'b0;
assign   tb_i_reset[488]                      =   1'b0;
assign   tb_i_sop[488]                        =   1'b0;
assign   tb_i_key_update[488]                 =   1'b0;
assign   tb_i_key[488]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[488]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[488]               =   1'b0;
assign   tb_i_rf_static_encrypt[488]          =   1'b1;
assign   tb_i_clear_fault_flags[488]          =   1'b0;
assign   tb_i_rf_static_aad_length[488]       =   64'h0000000000000100;
assign   tb_i_aad[488]                        =   tb_i_aad[487];
assign   tb_i_rf_static_plaintext_length[488] =   64'h0000000000000280;
assign   tb_i_plaintext[488]                  =   tb_i_plaintext[487];
assign   tb_o_valid[488]                      =   1'b0;
assign   tb_o_sop[488]                        =   1'b0;
assign   tb_o_ciphertext[488]                 =   tb_o_ciphertext[487];
assign   tb_o_tag_ready[488]                  =   1'b0;
assign   tb_o_tag[488]                        =   tb_o_tag[487];

// CLK no. 489/1240
// *************************************************
assign   tb_i_valid[489]                      =   1'b0;
assign   tb_i_reset[489]                      =   1'b0;
assign   tb_i_sop[489]                        =   1'b0;
assign   tb_i_key_update[489]                 =   1'b0;
assign   tb_i_key[489]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[489]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[489]               =   1'b0;
assign   tb_i_rf_static_encrypt[489]          =   1'b1;
assign   tb_i_clear_fault_flags[489]          =   1'b0;
assign   tb_i_rf_static_aad_length[489]       =   64'h0000000000000100;
assign   tb_i_aad[489]                        =   tb_i_aad[488];
assign   tb_i_rf_static_plaintext_length[489] =   64'h0000000000000280;
assign   tb_i_plaintext[489]                  =   tb_i_plaintext[488];
assign   tb_o_valid[489]                      =   1'b0;
assign   tb_o_sop[489]                        =   1'b0;
assign   tb_o_ciphertext[489]                 =   tb_o_ciphertext[488];
assign   tb_o_tag_ready[489]                  =   1'b0;
assign   tb_o_tag[489]                        =   tb_o_tag[488];

// CLK no. 490/1240
// *************************************************
assign   tb_i_valid[490]                      =   1'b0;
assign   tb_i_reset[490]                      =   1'b0;
assign   tb_i_sop[490]                        =   1'b0;
assign   tb_i_key_update[490]                 =   1'b0;
assign   tb_i_key[490]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[490]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[490]               =   1'b0;
assign   tb_i_rf_static_encrypt[490]          =   1'b1;
assign   tb_i_clear_fault_flags[490]          =   1'b0;
assign   tb_i_rf_static_aad_length[490]       =   64'h0000000000000100;
assign   tb_i_aad[490]                        =   tb_i_aad[489];
assign   tb_i_rf_static_plaintext_length[490] =   64'h0000000000000280;
assign   tb_i_plaintext[490]                  =   tb_i_plaintext[489];
assign   tb_o_valid[490]                      =   1'b0;
assign   tb_o_sop[490]                        =   1'b0;
assign   tb_o_ciphertext[490]                 =   tb_o_ciphertext[489];
assign   tb_o_tag_ready[490]                  =   1'b0;
assign   tb_o_tag[490]                        =   tb_o_tag[489];

// CLK no. 491/1240
// *************************************************
assign   tb_i_valid[491]                      =   1'b0;
assign   tb_i_reset[491]                      =   1'b0;
assign   tb_i_sop[491]                        =   1'b0;
assign   tb_i_key_update[491]                 =   1'b0;
assign   tb_i_key[491]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[491]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[491]               =   1'b0;
assign   tb_i_rf_static_encrypt[491]          =   1'b1;
assign   tb_i_clear_fault_flags[491]          =   1'b0;
assign   tb_i_rf_static_aad_length[491]       =   64'h0000000000000100;
assign   tb_i_aad[491]                        =   tb_i_aad[490];
assign   tb_i_rf_static_plaintext_length[491] =   64'h0000000000000280;
assign   tb_i_plaintext[491]                  =   tb_i_plaintext[490];
assign   tb_o_valid[491]                      =   1'b0;
assign   tb_o_sop[491]                        =   1'b0;
assign   tb_o_ciphertext[491]                 =   tb_o_ciphertext[490];
assign   tb_o_tag_ready[491]                  =   1'b0;
assign   tb_o_tag[491]                        =   tb_o_tag[490];

// CLK no. 492/1240
// *************************************************
assign   tb_i_valid[492]                      =   1'b0;
assign   tb_i_reset[492]                      =   1'b0;
assign   tb_i_sop[492]                        =   1'b0;
assign   tb_i_key_update[492]                 =   1'b0;
assign   tb_i_key[492]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[492]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[492]               =   1'b0;
assign   tb_i_rf_static_encrypt[492]          =   1'b1;
assign   tb_i_clear_fault_flags[492]          =   1'b0;
assign   tb_i_rf_static_aad_length[492]       =   64'h0000000000000100;
assign   tb_i_aad[492]                        =   tb_i_aad[491];
assign   tb_i_rf_static_plaintext_length[492] =   64'h0000000000000280;
assign   tb_i_plaintext[492]                  =   tb_i_plaintext[491];
assign   tb_o_valid[492]                      =   1'b0;
assign   tb_o_sop[492]                        =   1'b0;
assign   tb_o_ciphertext[492]                 =   tb_o_ciphertext[491];
assign   tb_o_tag_ready[492]                  =   1'b0;
assign   tb_o_tag[492]                        =   tb_o_tag[491];

// CLK no. 493/1240
// *************************************************
assign   tb_i_valid[493]                      =   1'b0;
assign   tb_i_reset[493]                      =   1'b0;
assign   tb_i_sop[493]                        =   1'b0;
assign   tb_i_key_update[493]                 =   1'b0;
assign   tb_i_key[493]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[493]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[493]               =   1'b0;
assign   tb_i_rf_static_encrypt[493]          =   1'b1;
assign   tb_i_clear_fault_flags[493]          =   1'b0;
assign   tb_i_rf_static_aad_length[493]       =   64'h0000000000000100;
assign   tb_i_aad[493]                        =   tb_i_aad[492];
assign   tb_i_rf_static_plaintext_length[493] =   64'h0000000000000280;
assign   tb_i_plaintext[493]                  =   tb_i_plaintext[492];
assign   tb_o_valid[493]                      =   1'b0;
assign   tb_o_sop[493]                        =   1'b0;
assign   tb_o_ciphertext[493]                 =   tb_o_ciphertext[492];
assign   tb_o_tag_ready[493]                  =   1'b0;
assign   tb_o_tag[493]                        =   tb_o_tag[492];

// CLK no. 494/1240
// *************************************************
assign   tb_i_valid[494]                      =   1'b0;
assign   tb_i_reset[494]                      =   1'b0;
assign   tb_i_sop[494]                        =   1'b0;
assign   tb_i_key_update[494]                 =   1'b0;
assign   tb_i_key[494]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[494]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[494]               =   1'b0;
assign   tb_i_rf_static_encrypt[494]          =   1'b1;
assign   tb_i_clear_fault_flags[494]          =   1'b0;
assign   tb_i_rf_static_aad_length[494]       =   64'h0000000000000100;
assign   tb_i_aad[494]                        =   tb_i_aad[493];
assign   tb_i_rf_static_plaintext_length[494] =   64'h0000000000000280;
assign   tb_i_plaintext[494]                  =   tb_i_plaintext[493];
assign   tb_o_valid[494]                      =   1'b0;
assign   tb_o_sop[494]                        =   1'b0;
assign   tb_o_ciphertext[494]                 =   tb_o_ciphertext[493];
assign   tb_o_tag_ready[494]                  =   1'b0;
assign   tb_o_tag[494]                        =   tb_o_tag[493];

// CLK no. 495/1240
// *************************************************
assign   tb_i_valid[495]                      =   1'b0;
assign   tb_i_reset[495]                      =   1'b0;
assign   tb_i_sop[495]                        =   1'b0;
assign   tb_i_key_update[495]                 =   1'b0;
assign   tb_i_key[495]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[495]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[495]               =   1'b0;
assign   tb_i_rf_static_encrypt[495]          =   1'b1;
assign   tb_i_clear_fault_flags[495]          =   1'b0;
assign   tb_i_rf_static_aad_length[495]       =   64'h0000000000000100;
assign   tb_i_aad[495]                        =   tb_i_aad[494];
assign   tb_i_rf_static_plaintext_length[495] =   64'h0000000000000280;
assign   tb_i_plaintext[495]                  =   tb_i_plaintext[494];
assign   tb_o_valid[495]                      =   1'b0;
assign   tb_o_sop[495]                        =   1'b0;
assign   tb_o_ciphertext[495]                 =   tb_o_ciphertext[494];
assign   tb_o_tag_ready[495]                  =   1'b0;
assign   tb_o_tag[495]                        =   tb_o_tag[494];

// CLK no. 496/1240
// *************************************************
assign   tb_i_valid[496]                      =   1'b0;
assign   tb_i_reset[496]                      =   1'b0;
assign   tb_i_sop[496]                        =   1'b0;
assign   tb_i_key_update[496]                 =   1'b0;
assign   tb_i_key[496]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[496]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[496]               =   1'b0;
assign   tb_i_rf_static_encrypt[496]          =   1'b1;
assign   tb_i_clear_fault_flags[496]          =   1'b0;
assign   tb_i_rf_static_aad_length[496]       =   64'h0000000000000100;
assign   tb_i_aad[496]                        =   tb_i_aad[495];
assign   tb_i_rf_static_plaintext_length[496] =   64'h0000000000000280;
assign   tb_i_plaintext[496]                  =   tb_i_plaintext[495];
assign   tb_o_valid[496]                      =   1'b0;
assign   tb_o_sop[496]                        =   1'b0;
assign   tb_o_ciphertext[496]                 =   tb_o_ciphertext[495];
assign   tb_o_tag_ready[496]                  =   1'b0;
assign   tb_o_tag[496]                        =   tb_o_tag[495];

// CLK no. 497/1240
// *************************************************
assign   tb_i_valid[497]                      =   1'b0;
assign   tb_i_reset[497]                      =   1'b0;
assign   tb_i_sop[497]                        =   1'b0;
assign   tb_i_key_update[497]                 =   1'b0;
assign   tb_i_key[497]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[497]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[497]               =   1'b0;
assign   tb_i_rf_static_encrypt[497]          =   1'b1;
assign   tb_i_clear_fault_flags[497]          =   1'b0;
assign   tb_i_rf_static_aad_length[497]       =   64'h0000000000000100;
assign   tb_i_aad[497]                        =   tb_i_aad[496];
assign   tb_i_rf_static_plaintext_length[497] =   64'h0000000000000280;
assign   tb_i_plaintext[497]                  =   tb_i_plaintext[496];
assign   tb_o_valid[497]                      =   1'b0;
assign   tb_o_sop[497]                        =   1'b0;
assign   tb_o_ciphertext[497]                 =   tb_o_ciphertext[496];
assign   tb_o_tag_ready[497]                  =   1'b0;
assign   tb_o_tag[497]                        =   tb_o_tag[496];

// CLK no. 498/1240
// *************************************************
assign   tb_i_valid[498]                      =   1'b0;
assign   tb_i_reset[498]                      =   1'b0;
assign   tb_i_sop[498]                        =   1'b0;
assign   tb_i_key_update[498]                 =   1'b0;
assign   tb_i_key[498]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[498]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[498]               =   1'b0;
assign   tb_i_rf_static_encrypt[498]          =   1'b1;
assign   tb_i_clear_fault_flags[498]          =   1'b0;
assign   tb_i_rf_static_aad_length[498]       =   64'h0000000000000100;
assign   tb_i_aad[498]                        =   tb_i_aad[497];
assign   tb_i_rf_static_plaintext_length[498] =   64'h0000000000000280;
assign   tb_i_plaintext[498]                  =   tb_i_plaintext[497];
assign   tb_o_valid[498]                      =   1'b0;
assign   tb_o_sop[498]                        =   1'b0;
assign   tb_o_ciphertext[498]                 =   tb_o_ciphertext[497];
assign   tb_o_tag_ready[498]                  =   1'b0;
assign   tb_o_tag[498]                        =   tb_o_tag[497];

// CLK no. 499/1240
// *************************************************
assign   tb_i_valid[499]                      =   1'b0;
assign   tb_i_reset[499]                      =   1'b0;
assign   tb_i_sop[499]                        =   1'b0;
assign   tb_i_key_update[499]                 =   1'b0;
assign   tb_i_key[499]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[499]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[499]               =   1'b0;
assign   tb_i_rf_static_encrypt[499]          =   1'b1;
assign   tb_i_clear_fault_flags[499]          =   1'b0;
assign   tb_i_rf_static_aad_length[499]       =   64'h0000000000000100;
assign   tb_i_aad[499]                        =   tb_i_aad[498];
assign   tb_i_rf_static_plaintext_length[499] =   64'h0000000000000280;
assign   tb_i_plaintext[499]                  =   tb_i_plaintext[498];
assign   tb_o_valid[499]                      =   1'b0;
assign   tb_o_sop[499]                        =   1'b0;
assign   tb_o_ciphertext[499]                 =   tb_o_ciphertext[498];
assign   tb_o_tag_ready[499]                  =   1'b0;
assign   tb_o_tag[499]                        =   tb_o_tag[498];

// CLK no. 500/1240
// *************************************************
assign   tb_i_valid[500]                      =   1'b0;
assign   tb_i_reset[500]                      =   1'b0;
assign   tb_i_sop[500]                        =   1'b0;
assign   tb_i_key_update[500]                 =   1'b0;
assign   tb_i_key[500]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[500]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[500]               =   1'b0;
assign   tb_i_rf_static_encrypt[500]          =   1'b1;
assign   tb_i_clear_fault_flags[500]          =   1'b0;
assign   tb_i_rf_static_aad_length[500]       =   64'h0000000000000100;
assign   tb_i_aad[500]                        =   tb_i_aad[499];
assign   tb_i_rf_static_plaintext_length[500] =   64'h0000000000000280;
assign   tb_i_plaintext[500]                  =   tb_i_plaintext[499];
assign   tb_o_valid[500]                      =   1'b0;
assign   tb_o_sop[500]                        =   1'b0;
assign   tb_o_ciphertext[500]                 =   tb_o_ciphertext[499];
assign   tb_o_tag_ready[500]                  =   1'b0;
assign   tb_o_tag[500]                        =   tb_o_tag[499];

// CLK no. 501/1240
// *************************************************
assign   tb_i_valid[501]                      =   1'b0;
assign   tb_i_reset[501]                      =   1'b0;
assign   tb_i_sop[501]                        =   1'b0;
assign   tb_i_key_update[501]                 =   1'b0;
assign   tb_i_key[501]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[501]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[501]               =   1'b0;
assign   tb_i_rf_static_encrypt[501]          =   1'b1;
assign   tb_i_clear_fault_flags[501]          =   1'b0;
assign   tb_i_rf_static_aad_length[501]       =   64'h0000000000000100;
assign   tb_i_aad[501]                        =   tb_i_aad[500];
assign   tb_i_rf_static_plaintext_length[501] =   64'h0000000000000280;
assign   tb_i_plaintext[501]                  =   tb_i_plaintext[500];
assign   tb_o_valid[501]                      =   1'b0;
assign   tb_o_sop[501]                        =   1'b0;
assign   tb_o_ciphertext[501]                 =   tb_o_ciphertext[500];
assign   tb_o_tag_ready[501]                  =   1'b0;
assign   tb_o_tag[501]                        =   tb_o_tag[500];

// CLK no. 502/1240
// *************************************************
assign   tb_i_valid[502]                      =   1'b0;
assign   tb_i_reset[502]                      =   1'b0;
assign   tb_i_sop[502]                        =   1'b0;
assign   tb_i_key_update[502]                 =   1'b0;
assign   tb_i_key[502]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[502]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[502]               =   1'b0;
assign   tb_i_rf_static_encrypt[502]          =   1'b1;
assign   tb_i_clear_fault_flags[502]          =   1'b0;
assign   tb_i_rf_static_aad_length[502]       =   64'h0000000000000100;
assign   tb_i_aad[502]                        =   tb_i_aad[501];
assign   tb_i_rf_static_plaintext_length[502] =   64'h0000000000000280;
assign   tb_i_plaintext[502]                  =   tb_i_plaintext[501];
assign   tb_o_valid[502]                      =   1'b0;
assign   tb_o_sop[502]                        =   1'b0;
assign   tb_o_ciphertext[502]                 =   tb_o_ciphertext[501];
assign   tb_o_tag_ready[502]                  =   1'b0;
assign   tb_o_tag[502]                        =   tb_o_tag[501];

// CLK no. 503/1240
// *************************************************
assign   tb_i_valid[503]                      =   1'b0;
assign   tb_i_reset[503]                      =   1'b0;
assign   tb_i_sop[503]                        =   1'b0;
assign   tb_i_key_update[503]                 =   1'b0;
assign   tb_i_key[503]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[503]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[503]               =   1'b0;
assign   tb_i_rf_static_encrypt[503]          =   1'b1;
assign   tb_i_clear_fault_flags[503]          =   1'b0;
assign   tb_i_rf_static_aad_length[503]       =   64'h0000000000000100;
assign   tb_i_aad[503]                        =   tb_i_aad[502];
assign   tb_i_rf_static_plaintext_length[503] =   64'h0000000000000280;
assign   tb_i_plaintext[503]                  =   tb_i_plaintext[502];
assign   tb_o_valid[503]                      =   1'b0;
assign   tb_o_sop[503]                        =   1'b0;
assign   tb_o_ciphertext[503]                 =   tb_o_ciphertext[502];
assign   tb_o_tag_ready[503]                  =   1'b0;
assign   tb_o_tag[503]                        =   tb_o_tag[502];

// CLK no. 504/1240
// *************************************************
assign   tb_i_valid[504]                      =   1'b0;
assign   tb_i_reset[504]                      =   1'b0;
assign   tb_i_sop[504]                        =   1'b0;
assign   tb_i_key_update[504]                 =   1'b0;
assign   tb_i_key[504]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[504]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[504]               =   1'b0;
assign   tb_i_rf_static_encrypt[504]          =   1'b1;
assign   tb_i_clear_fault_flags[504]          =   1'b0;
assign   tb_i_rf_static_aad_length[504]       =   64'h0000000000000100;
assign   tb_i_aad[504]                        =   tb_i_aad[503];
assign   tb_i_rf_static_plaintext_length[504] =   64'h0000000000000280;
assign   tb_i_plaintext[504]                  =   tb_i_plaintext[503];
assign   tb_o_valid[504]                      =   1'b0;
assign   tb_o_sop[504]                        =   1'b0;
assign   tb_o_ciphertext[504]                 =   tb_o_ciphertext[503];
assign   tb_o_tag_ready[504]                  =   1'b0;
assign   tb_o_tag[504]                        =   tb_o_tag[503];

// CLK no. 505/1240
// *************************************************
assign   tb_i_valid[505]                      =   1'b0;
assign   tb_i_reset[505]                      =   1'b0;
assign   tb_i_sop[505]                        =   1'b0;
assign   tb_i_key_update[505]                 =   1'b0;
assign   tb_i_key[505]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[505]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[505]               =   1'b0;
assign   tb_i_rf_static_encrypt[505]          =   1'b1;
assign   tb_i_clear_fault_flags[505]          =   1'b0;
assign   tb_i_rf_static_aad_length[505]       =   64'h0000000000000100;
assign   tb_i_aad[505]                        =   tb_i_aad[504];
assign   tb_i_rf_static_plaintext_length[505] =   64'h0000000000000280;
assign   tb_i_plaintext[505]                  =   tb_i_plaintext[504];
assign   tb_o_valid[505]                      =   1'b0;
assign   tb_o_sop[505]                        =   1'b0;
assign   tb_o_ciphertext[505]                 =   tb_o_ciphertext[504];
assign   tb_o_tag_ready[505]                  =   1'b0;
assign   tb_o_tag[505]                        =   tb_o_tag[504];

// CLK no. 506/1240
// *************************************************
assign   tb_i_valid[506]                      =   1'b0;
assign   tb_i_reset[506]                      =   1'b0;
assign   tb_i_sop[506]                        =   1'b0;
assign   tb_i_key_update[506]                 =   1'b0;
assign   tb_i_key[506]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[506]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[506]               =   1'b0;
assign   tb_i_rf_static_encrypt[506]          =   1'b1;
assign   tb_i_clear_fault_flags[506]          =   1'b0;
assign   tb_i_rf_static_aad_length[506]       =   64'h0000000000000100;
assign   tb_i_aad[506]                        =   tb_i_aad[505];
assign   tb_i_rf_static_plaintext_length[506] =   64'h0000000000000280;
assign   tb_i_plaintext[506]                  =   tb_i_plaintext[505];
assign   tb_o_valid[506]                      =   1'b0;
assign   tb_o_sop[506]                        =   1'b0;
assign   tb_o_ciphertext[506]                 =   tb_o_ciphertext[505];
assign   tb_o_tag_ready[506]                  =   1'b0;
assign   tb_o_tag[506]                        =   tb_o_tag[505];

// CLK no. 507/1240
// *************************************************
assign   tb_i_valid[507]                      =   1'b0;
assign   tb_i_reset[507]                      =   1'b0;
assign   tb_i_sop[507]                        =   1'b0;
assign   tb_i_key_update[507]                 =   1'b0;
assign   tb_i_key[507]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[507]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[507]               =   1'b0;
assign   tb_i_rf_static_encrypt[507]          =   1'b1;
assign   tb_i_clear_fault_flags[507]          =   1'b0;
assign   tb_i_rf_static_aad_length[507]       =   64'h0000000000000100;
assign   tb_i_aad[507]                        =   tb_i_aad[506];
assign   tb_i_rf_static_plaintext_length[507] =   64'h0000000000000280;
assign   tb_i_plaintext[507]                  =   tb_i_plaintext[506];
assign   tb_o_valid[507]                      =   1'b0;
assign   tb_o_sop[507]                        =   1'b0;
assign   tb_o_ciphertext[507]                 =   tb_o_ciphertext[506];
assign   tb_o_tag_ready[507]                  =   1'b0;
assign   tb_o_tag[507]                        =   tb_o_tag[506];

// CLK no. 508/1240
// *************************************************
assign   tb_i_valid[508]                      =   1'b0;
assign   tb_i_reset[508]                      =   1'b0;
assign   tb_i_sop[508]                        =   1'b0;
assign   tb_i_key_update[508]                 =   1'b0;
assign   tb_i_key[508]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[508]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[508]               =   1'b0;
assign   tb_i_rf_static_encrypt[508]          =   1'b1;
assign   tb_i_clear_fault_flags[508]          =   1'b0;
assign   tb_i_rf_static_aad_length[508]       =   64'h0000000000000100;
assign   tb_i_aad[508]                        =   tb_i_aad[507];
assign   tb_i_rf_static_plaintext_length[508] =   64'h0000000000000280;
assign   tb_i_plaintext[508]                  =   tb_i_plaintext[507];
assign   tb_o_valid[508]                      =   1'b0;
assign   tb_o_sop[508]                        =   1'b0;
assign   tb_o_ciphertext[508]                 =   tb_o_ciphertext[507];
assign   tb_o_tag_ready[508]                  =   1'b0;
assign   tb_o_tag[508]                        =   tb_o_tag[507];

// CLK no. 509/1240
// *************************************************
assign   tb_i_valid[509]                      =   1'b0;
assign   tb_i_reset[509]                      =   1'b0;
assign   tb_i_sop[509]                        =   1'b0;
assign   tb_i_key_update[509]                 =   1'b0;
assign   tb_i_key[509]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[509]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[509]               =   1'b0;
assign   tb_i_rf_static_encrypt[509]          =   1'b1;
assign   tb_i_clear_fault_flags[509]          =   1'b0;
assign   tb_i_rf_static_aad_length[509]       =   64'h0000000000000100;
assign   tb_i_aad[509]                        =   tb_i_aad[508];
assign   tb_i_rf_static_plaintext_length[509] =   64'h0000000000000280;
assign   tb_i_plaintext[509]                  =   tb_i_plaintext[508];
assign   tb_o_valid[509]                      =   1'b0;
assign   tb_o_sop[509]                        =   1'b0;
assign   tb_o_ciphertext[509]                 =   tb_o_ciphertext[508];
assign   tb_o_tag_ready[509]                  =   1'b0;
assign   tb_o_tag[509]                        =   tb_o_tag[508];

// CLK no. 510/1240
// *************************************************
assign   tb_i_valid[510]                      =   1'b0;
assign   tb_i_reset[510]                      =   1'b0;
assign   tb_i_sop[510]                        =   1'b0;
assign   tb_i_key_update[510]                 =   1'b0;
assign   tb_i_key[510]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[510]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[510]               =   1'b0;
assign   tb_i_rf_static_encrypt[510]          =   1'b1;
assign   tb_i_clear_fault_flags[510]          =   1'b0;
assign   tb_i_rf_static_aad_length[510]       =   64'h0000000000000100;
assign   tb_i_aad[510]                        =   tb_i_aad[509];
assign   tb_i_rf_static_plaintext_length[510] =   64'h0000000000000280;
assign   tb_i_plaintext[510]                  =   tb_i_plaintext[509];
assign   tb_o_valid[510]                      =   1'b0;
assign   tb_o_sop[510]                        =   1'b0;
assign   tb_o_ciphertext[510]                 =   tb_o_ciphertext[509];
assign   tb_o_tag_ready[510]                  =   1'b0;
assign   tb_o_tag[510]                        =   tb_o_tag[509];

// CLK no. 511/1240
// *************************************************
assign   tb_i_valid[511]                      =   1'b0;
assign   tb_i_reset[511]                      =   1'b0;
assign   tb_i_sop[511]                        =   1'b0;
assign   tb_i_key_update[511]                 =   1'b0;
assign   tb_i_key[511]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[511]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[511]               =   1'b0;
assign   tb_i_rf_static_encrypt[511]          =   1'b1;
assign   tb_i_clear_fault_flags[511]          =   1'b0;
assign   tb_i_rf_static_aad_length[511]       =   64'h0000000000000100;
assign   tb_i_aad[511]                        =   tb_i_aad[510];
assign   tb_i_rf_static_plaintext_length[511] =   64'h0000000000000280;
assign   tb_i_plaintext[511]                  =   tb_i_plaintext[510];
assign   tb_o_valid[511]                      =   1'b0;
assign   tb_o_sop[511]                        =   1'b0;
assign   tb_o_ciphertext[511]                 =   tb_o_ciphertext[510];
assign   tb_o_tag_ready[511]                  =   1'b0;
assign   tb_o_tag[511]                        =   tb_o_tag[510];

// CLK no. 512/1240
// *************************************************
assign   tb_i_valid[512]                      =   1'b0;
assign   tb_i_reset[512]                      =   1'b0;
assign   tb_i_sop[512]                        =   1'b0;
assign   tb_i_key_update[512]                 =   1'b0;
assign   tb_i_key[512]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[512]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[512]               =   1'b0;
assign   tb_i_rf_static_encrypt[512]          =   1'b1;
assign   tb_i_clear_fault_flags[512]          =   1'b0;
assign   tb_i_rf_static_aad_length[512]       =   64'h0000000000000100;
assign   tb_i_aad[512]                        =   tb_i_aad[511];
assign   tb_i_rf_static_plaintext_length[512] =   64'h0000000000000280;
assign   tb_i_plaintext[512]                  =   tb_i_plaintext[511];
assign   tb_o_valid[512]                      =   1'b0;
assign   tb_o_sop[512]                        =   1'b0;
assign   tb_o_ciphertext[512]                 =   tb_o_ciphertext[511];
assign   tb_o_tag_ready[512]                  =   1'b0;
assign   tb_o_tag[512]                        =   tb_o_tag[511];

// CLK no. 513/1240
// *************************************************
assign   tb_i_valid[513]                      =   1'b0;
assign   tb_i_reset[513]                      =   1'b0;
assign   tb_i_sop[513]                        =   1'b0;
assign   tb_i_key_update[513]                 =   1'b0;
assign   tb_i_key[513]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[513]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[513]               =   1'b0;
assign   tb_i_rf_static_encrypt[513]          =   1'b1;
assign   tb_i_clear_fault_flags[513]          =   1'b0;
assign   tb_i_rf_static_aad_length[513]       =   64'h0000000000000100;
assign   tb_i_aad[513]                        =   tb_i_aad[512];
assign   tb_i_rf_static_plaintext_length[513] =   64'h0000000000000280;
assign   tb_i_plaintext[513]                  =   tb_i_plaintext[512];
assign   tb_o_valid[513]                      =   1'b0;
assign   tb_o_sop[513]                        =   1'b0;
assign   tb_o_ciphertext[513]                 =   tb_o_ciphertext[512];
assign   tb_o_tag_ready[513]                  =   1'b0;
assign   tb_o_tag[513]                        =   tb_o_tag[512];

// CLK no. 514/1240
// *************************************************
assign   tb_i_valid[514]                      =   1'b0;
assign   tb_i_reset[514]                      =   1'b0;
assign   tb_i_sop[514]                        =   1'b0;
assign   tb_i_key_update[514]                 =   1'b0;
assign   tb_i_key[514]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[514]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[514]               =   1'b0;
assign   tb_i_rf_static_encrypt[514]          =   1'b1;
assign   tb_i_clear_fault_flags[514]          =   1'b0;
assign   tb_i_rf_static_aad_length[514]       =   64'h0000000000000100;
assign   tb_i_aad[514]                        =   tb_i_aad[513];
assign   tb_i_rf_static_plaintext_length[514] =   64'h0000000000000280;
assign   tb_i_plaintext[514]                  =   tb_i_plaintext[513];
assign   tb_o_valid[514]                      =   1'b0;
assign   tb_o_sop[514]                        =   1'b0;
assign   tb_o_ciphertext[514]                 =   tb_o_ciphertext[513];
assign   tb_o_tag_ready[514]                  =   1'b0;
assign   tb_o_tag[514]                        =   tb_o_tag[513];

// CLK no. 515/1240
// *************************************************
assign   tb_i_valid[515]                      =   1'b0;
assign   tb_i_reset[515]                      =   1'b0;
assign   tb_i_sop[515]                        =   1'b0;
assign   tb_i_key_update[515]                 =   1'b0;
assign   tb_i_key[515]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[515]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[515]               =   1'b0;
assign   tb_i_rf_static_encrypt[515]          =   1'b1;
assign   tb_i_clear_fault_flags[515]          =   1'b0;
assign   tb_i_rf_static_aad_length[515]       =   64'h0000000000000100;
assign   tb_i_aad[515]                        =   tb_i_aad[514];
assign   tb_i_rf_static_plaintext_length[515] =   64'h0000000000000280;
assign   tb_i_plaintext[515]                  =   tb_i_plaintext[514];
assign   tb_o_valid[515]                      =   1'b0;
assign   tb_o_sop[515]                        =   1'b0;
assign   tb_o_ciphertext[515]                 =   tb_o_ciphertext[514];
assign   tb_o_tag_ready[515]                  =   1'b0;
assign   tb_o_tag[515]                        =   tb_o_tag[514];

// CLK no. 516/1240
// *************************************************
assign   tb_i_valid[516]                      =   1'b0;
assign   tb_i_reset[516]                      =   1'b0;
assign   tb_i_sop[516]                        =   1'b0;
assign   tb_i_key_update[516]                 =   1'b0;
assign   tb_i_key[516]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[516]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[516]               =   1'b0;
assign   tb_i_rf_static_encrypt[516]          =   1'b1;
assign   tb_i_clear_fault_flags[516]          =   1'b0;
assign   tb_i_rf_static_aad_length[516]       =   64'h0000000000000100;
assign   tb_i_aad[516]                        =   tb_i_aad[515];
assign   tb_i_rf_static_plaintext_length[516] =   64'h0000000000000280;
assign   tb_i_plaintext[516]                  =   tb_i_plaintext[515];
assign   tb_o_valid[516]                      =   1'b0;
assign   tb_o_sop[516]                        =   1'b0;
assign   tb_o_ciphertext[516]                 =   tb_o_ciphertext[515];
assign   tb_o_tag_ready[516]                  =   1'b0;
assign   tb_o_tag[516]                        =   tb_o_tag[515];

// CLK no. 517/1240
// *************************************************
assign   tb_i_valid[517]                      =   1'b0;
assign   tb_i_reset[517]                      =   1'b0;
assign   tb_i_sop[517]                        =   1'b0;
assign   tb_i_key_update[517]                 =   1'b0;
assign   tb_i_key[517]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[517]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[517]               =   1'b0;
assign   tb_i_rf_static_encrypt[517]          =   1'b1;
assign   tb_i_clear_fault_flags[517]          =   1'b0;
assign   tb_i_rf_static_aad_length[517]       =   64'h0000000000000100;
assign   tb_i_aad[517]                        =   tb_i_aad[516];
assign   tb_i_rf_static_plaintext_length[517] =   64'h0000000000000280;
assign   tb_i_plaintext[517]                  =   tb_i_plaintext[516];
assign   tb_o_valid[517]                      =   1'b0;
assign   tb_o_sop[517]                        =   1'b0;
assign   tb_o_ciphertext[517]                 =   tb_o_ciphertext[516];
assign   tb_o_tag_ready[517]                  =   1'b0;
assign   tb_o_tag[517]                        =   tb_o_tag[516];

// CLK no. 518/1240
// *************************************************
assign   tb_i_valid[518]                      =   1'b0;
assign   tb_i_reset[518]                      =   1'b0;
assign   tb_i_sop[518]                        =   1'b0;
assign   tb_i_key_update[518]                 =   1'b0;
assign   tb_i_key[518]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[518]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[518]               =   1'b0;
assign   tb_i_rf_static_encrypt[518]          =   1'b1;
assign   tb_i_clear_fault_flags[518]          =   1'b0;
assign   tb_i_rf_static_aad_length[518]       =   64'h0000000000000100;
assign   tb_i_aad[518]                        =   tb_i_aad[517];
assign   tb_i_rf_static_plaintext_length[518] =   64'h0000000000000280;
assign   tb_i_plaintext[518]                  =   tb_i_plaintext[517];
assign   tb_o_valid[518]                      =   1'b0;
assign   tb_o_sop[518]                        =   1'b0;
assign   tb_o_ciphertext[518]                 =   tb_o_ciphertext[517];
assign   tb_o_tag_ready[518]                  =   1'b0;
assign   tb_o_tag[518]                        =   tb_o_tag[517];

// CLK no. 519/1240
// *************************************************
assign   tb_i_valid[519]                      =   1'b0;
assign   tb_i_reset[519]                      =   1'b0;
assign   tb_i_sop[519]                        =   1'b0;
assign   tb_i_key_update[519]                 =   1'b0;
assign   tb_i_key[519]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[519]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[519]               =   1'b0;
assign   tb_i_rf_static_encrypt[519]          =   1'b1;
assign   tb_i_clear_fault_flags[519]          =   1'b0;
assign   tb_i_rf_static_aad_length[519]       =   64'h0000000000000100;
assign   tb_i_aad[519]                        =   tb_i_aad[518];
assign   tb_i_rf_static_plaintext_length[519] =   64'h0000000000000280;
assign   tb_i_plaintext[519]                  =   tb_i_plaintext[518];
assign   tb_o_valid[519]                      =   1'b1;
assign   tb_o_sop[519]                        =   1'b1;
assign   tb_o_ciphertext[519]                 =   256'h7864ade9957f67eb9a88e2a668ca97f5b16276dfd75ae81a1e96b92f8969d7df;
assign   tb_o_tag_ready[519]                  =   1'b0;
assign   tb_o_tag[519]                        =   tb_o_tag[518];

// CLK no. 520/1240
// *************************************************
assign   tb_i_valid[520]                      =   1'b0;
assign   tb_i_reset[520]                      =   1'b0;
assign   tb_i_sop[520]                        =   1'b0;
assign   tb_i_key_update[520]                 =   1'b0;
assign   tb_i_key[520]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[520]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[520]               =   1'b0;
assign   tb_i_rf_static_encrypt[520]          =   1'b1;
assign   tb_i_clear_fault_flags[520]          =   1'b0;
assign   tb_i_rf_static_aad_length[520]       =   64'h0000000000000100;
assign   tb_i_aad[520]                        =   tb_i_aad[519];
assign   tb_i_rf_static_plaintext_length[520] =   64'h0000000000000280;
assign   tb_i_plaintext[520]                  =   tb_i_plaintext[519];
assign   tb_o_valid[520]                      =   1'b1;
assign   tb_o_sop[520]                        =   1'b0;
assign   tb_o_ciphertext[520]                 =   256'h7eb12f642d3c1abcaf93e2b5fe7aaf0f099a9e25083a9c849f65b1e69e6d098b;
assign   tb_o_tag_ready[520]                  =   1'b0;
assign   tb_o_tag[520]                        =   tb_o_tag[519];

// CLK no. 521/1240
// *************************************************
assign   tb_i_valid[521]                      =   1'b0;
assign   tb_i_reset[521]                      =   1'b0;
assign   tb_i_sop[521]                        =   1'b0;
assign   tb_i_key_update[521]                 =   1'b0;
assign   tb_i_key[521]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[521]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[521]               =   1'b0;
assign   tb_i_rf_static_encrypt[521]          =   1'b1;
assign   tb_i_clear_fault_flags[521]          =   1'b0;
assign   tb_i_rf_static_aad_length[521]       =   64'h0000000000000100;
assign   tb_i_aad[521]                        =   tb_i_aad[520];
assign   tb_i_rf_static_plaintext_length[521] =   64'h0000000000000280;
assign   tb_i_plaintext[521]                  =   tb_i_plaintext[520];
assign   tb_o_valid[521]                      =   1'b1;
assign   tb_o_sop[521]                        =   1'b0;
assign   tb_o_ciphertext[521]                 =   256'hc201fb7b847285eb7d9db9dffff337a5;
assign   tb_o_tag_ready[521]                  =   1'b0;
assign   tb_o_tag[521]                        =   tb_o_tag[520];

// CLK no. 522/1240
// *************************************************
assign   tb_i_valid[522]                      =   1'b0;
assign   tb_i_reset[522]                      =   1'b0;
assign   tb_i_sop[522]                        =   1'b0;
assign   tb_i_key_update[522]                 =   1'b0;
assign   tb_i_key[522]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[522]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[522]               =   1'b0;
assign   tb_i_rf_static_encrypt[522]          =   1'b1;
assign   tb_i_clear_fault_flags[522]          =   1'b0;
assign   tb_i_rf_static_aad_length[522]       =   64'h0000000000000100;
assign   tb_i_aad[522]                        =   tb_i_aad[521];
assign   tb_i_rf_static_plaintext_length[522] =   64'h0000000000000280;
assign   tb_i_plaintext[522]                  =   tb_i_plaintext[521];
assign   tb_o_valid[522]                      =   1'b0;
assign   tb_o_sop[522]                        =   1'b0;
assign   tb_o_ciphertext[522]                 =   tb_o_ciphertext[521];
assign   tb_o_tag_ready[522]                  =   1'b0;
assign   tb_o_tag[522]                        =   tb_o_tag[521];

// CLK no. 523/1240
// *************************************************
assign   tb_i_valid[523]                      =   1'b0;
assign   tb_i_reset[523]                      =   1'b0;
assign   tb_i_sop[523]                        =   1'b0;
assign   tb_i_key_update[523]                 =   1'b0;
assign   tb_i_key[523]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[523]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[523]               =   1'b0;
assign   tb_i_rf_static_encrypt[523]          =   1'b1;
assign   tb_i_clear_fault_flags[523]          =   1'b0;
assign   tb_i_rf_static_aad_length[523]       =   64'h0000000000000100;
assign   tb_i_aad[523]                        =   tb_i_aad[522];
assign   tb_i_rf_static_plaintext_length[523] =   64'h0000000000000280;
assign   tb_i_plaintext[523]                  =   tb_i_plaintext[522];
assign   tb_o_valid[523]                      =   1'b0;
assign   tb_o_sop[523]                        =   1'b0;
assign   tb_o_ciphertext[523]                 =   tb_o_ciphertext[522];
assign   tb_o_tag_ready[523]                  =   1'b0;
assign   tb_o_tag[523]                        =   tb_o_tag[522];

// CLK no. 524/1240
// *************************************************
assign   tb_i_valid[524]                      =   1'b0;
assign   tb_i_reset[524]                      =   1'b0;
assign   tb_i_sop[524]                        =   1'b0;
assign   tb_i_key_update[524]                 =   1'b0;
assign   tb_i_key[524]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[524]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[524]               =   1'b0;
assign   tb_i_rf_static_encrypt[524]          =   1'b1;
assign   tb_i_clear_fault_flags[524]          =   1'b0;
assign   tb_i_rf_static_aad_length[524]       =   64'h0000000000000100;
assign   tb_i_aad[524]                        =   tb_i_aad[523];
assign   tb_i_rf_static_plaintext_length[524] =   64'h0000000000000280;
assign   tb_i_plaintext[524]                  =   tb_i_plaintext[523];
assign   tb_o_valid[524]                      =   1'b0;
assign   tb_o_sop[524]                        =   1'b0;
assign   tb_o_ciphertext[524]                 =   tb_o_ciphertext[523];
assign   tb_o_tag_ready[524]                  =   1'b0;
assign   tb_o_tag[524]                        =   tb_o_tag[523];

// CLK no. 525/1240
// *************************************************
assign   tb_i_valid[525]                      =   1'b0;
assign   tb_i_reset[525]                      =   1'b0;
assign   tb_i_sop[525]                        =   1'b0;
assign   tb_i_key_update[525]                 =   1'b0;
assign   tb_i_key[525]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[525]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[525]               =   1'b0;
assign   tb_i_rf_static_encrypt[525]          =   1'b1;
assign   tb_i_clear_fault_flags[525]          =   1'b0;
assign   tb_i_rf_static_aad_length[525]       =   64'h0000000000000100;
assign   tb_i_aad[525]                        =   tb_i_aad[524];
assign   tb_i_rf_static_plaintext_length[525] =   64'h0000000000000280;
assign   tb_i_plaintext[525]                  =   tb_i_plaintext[524];
assign   tb_o_valid[525]                      =   1'b0;
assign   tb_o_sop[525]                        =   1'b0;
assign   tb_o_ciphertext[525]                 =   tb_o_ciphertext[524];
assign   tb_o_tag_ready[525]                  =   1'b0;
assign   tb_o_tag[525]                        =   tb_o_tag[524];

// CLK no. 526/1240
// *************************************************
assign   tb_i_valid[526]                      =   1'b0;
assign   tb_i_reset[526]                      =   1'b0;
assign   tb_i_sop[526]                        =   1'b0;
assign   tb_i_key_update[526]                 =   1'b0;
assign   tb_i_key[526]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[526]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[526]               =   1'b0;
assign   tb_i_rf_static_encrypt[526]          =   1'b1;
assign   tb_i_clear_fault_flags[526]          =   1'b0;
assign   tb_i_rf_static_aad_length[526]       =   64'h0000000000000100;
assign   tb_i_aad[526]                        =   tb_i_aad[525];
assign   tb_i_rf_static_plaintext_length[526] =   64'h0000000000000280;
assign   tb_i_plaintext[526]                  =   tb_i_plaintext[525];
assign   tb_o_valid[526]                      =   1'b0;
assign   tb_o_sop[526]                        =   1'b0;
assign   tb_o_ciphertext[526]                 =   tb_o_ciphertext[525];
assign   tb_o_tag_ready[526]                  =   1'b0;
assign   tb_o_tag[526]                        =   tb_o_tag[525];

// CLK no. 527/1240
// *************************************************
assign   tb_i_valid[527]                      =   1'b0;
assign   tb_i_reset[527]                      =   1'b0;
assign   tb_i_sop[527]                        =   1'b0;
assign   tb_i_key_update[527]                 =   1'b0;
assign   tb_i_key[527]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[527]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[527]               =   1'b0;
assign   tb_i_rf_static_encrypt[527]          =   1'b1;
assign   tb_i_clear_fault_flags[527]          =   1'b0;
assign   tb_i_rf_static_aad_length[527]       =   64'h0000000000000100;
assign   tb_i_aad[527]                        =   tb_i_aad[526];
assign   tb_i_rf_static_plaintext_length[527] =   64'h0000000000000280;
assign   tb_i_plaintext[527]                  =   tb_i_plaintext[526];
assign   tb_o_valid[527]                      =   1'b0;
assign   tb_o_sop[527]                        =   1'b0;
assign   tb_o_ciphertext[527]                 =   tb_o_ciphertext[526];
assign   tb_o_tag_ready[527]                  =   1'b0;
assign   tb_o_tag[527]                        =   tb_o_tag[526];

// CLK no. 528/1240
// *************************************************
assign   tb_i_valid[528]                      =   1'b0;
assign   tb_i_reset[528]                      =   1'b0;
assign   tb_i_sop[528]                        =   1'b0;
assign   tb_i_key_update[528]                 =   1'b0;
assign   tb_i_key[528]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[528]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[528]               =   1'b0;
assign   tb_i_rf_static_encrypt[528]          =   1'b1;
assign   tb_i_clear_fault_flags[528]          =   1'b0;
assign   tb_i_rf_static_aad_length[528]       =   64'h0000000000000100;
assign   tb_i_aad[528]                        =   tb_i_aad[527];
assign   tb_i_rf_static_plaintext_length[528] =   64'h0000000000000280;
assign   tb_i_plaintext[528]                  =   tb_i_plaintext[527];
assign   tb_o_valid[528]                      =   1'b0;
assign   tb_o_sop[528]                        =   1'b0;
assign   tb_o_ciphertext[528]                 =   tb_o_ciphertext[527];
assign   tb_o_tag_ready[528]                  =   1'b0;
assign   tb_o_tag[528]                        =   tb_o_tag[527];

// CLK no. 529/1240
// *************************************************
assign   tb_i_valid[529]                      =   1'b0;
assign   tb_i_reset[529]                      =   1'b0;
assign   tb_i_sop[529]                        =   1'b0;
assign   tb_i_key_update[529]                 =   1'b0;
assign   tb_i_key[529]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[529]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[529]               =   1'b0;
assign   tb_i_rf_static_encrypt[529]          =   1'b1;
assign   tb_i_clear_fault_flags[529]          =   1'b0;
assign   tb_i_rf_static_aad_length[529]       =   64'h0000000000000100;
assign   tb_i_aad[529]                        =   tb_i_aad[528];
assign   tb_i_rf_static_plaintext_length[529] =   64'h0000000000000280;
assign   tb_i_plaintext[529]                  =   tb_i_plaintext[528];
assign   tb_o_valid[529]                      =   1'b0;
assign   tb_o_sop[529]                        =   1'b0;
assign   tb_o_ciphertext[529]                 =   tb_o_ciphertext[528];
assign   tb_o_tag_ready[529]                  =   1'b1;
assign   tb_o_tag[529]                        =   128'hccbb1712f6e0c2256c08577a38d462dc;

// CLK no. 530/1240
// *************************************************
assign   tb_i_valid[530]                      =   1'b0;
assign   tb_i_reset[530]                      =   1'b0;
assign   tb_i_sop[530]                        =   1'b0;
assign   tb_i_key_update[530]                 =   1'b0;
assign   tb_i_key[530]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[530]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[530]               =   1'b0;
assign   tb_i_rf_static_encrypt[530]          =   1'b1;
assign   tb_i_clear_fault_flags[530]          =   1'b0;
assign   tb_i_rf_static_aad_length[530]       =   64'h0000000000000100;
assign   tb_i_aad[530]                        =   tb_i_aad[529];
assign   tb_i_rf_static_plaintext_length[530] =   64'h0000000000000280;
assign   tb_i_plaintext[530]                  =   tb_i_plaintext[529];
assign   tb_o_valid[530]                      =   1'b0;
assign   tb_o_sop[530]                        =   1'b0;
assign   tb_o_ciphertext[530]                 =   tb_o_ciphertext[529];
assign   tb_o_tag_ready[530]                  =   1'b0;
assign   tb_o_tag[530]                        =   tb_o_tag[529];

// CLK no. 531/1240
// *************************************************
assign   tb_i_valid[531]                      =   1'b0;
assign   tb_i_reset[531]                      =   1'b0;
assign   tb_i_sop[531]                        =   1'b0;
assign   tb_i_key_update[531]                 =   1'b0;
assign   tb_i_key[531]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[531]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[531]               =   1'b0;
assign   tb_i_rf_static_encrypt[531]          =   1'b1;
assign   tb_i_clear_fault_flags[531]          =   1'b0;
assign   tb_i_rf_static_aad_length[531]       =   64'h0000000000000100;
assign   tb_i_aad[531]                        =   tb_i_aad[530];
assign   tb_i_rf_static_plaintext_length[531] =   64'h0000000000000280;
assign   tb_i_plaintext[531]                  =   tb_i_plaintext[530];
assign   tb_o_valid[531]                      =   1'b0;
assign   tb_o_sop[531]                        =   1'b0;
assign   tb_o_ciphertext[531]                 =   tb_o_ciphertext[530];
assign   tb_o_tag_ready[531]                  =   1'b0;
assign   tb_o_tag[531]                        =   tb_o_tag[530];

// CLK no. 532/1240
// *************************************************
assign   tb_i_valid[532]                      =   1'b0;
assign   tb_i_reset[532]                      =   1'b0;
assign   tb_i_sop[532]                        =   1'b1;
assign   tb_i_key_update[532]                 =   1'b0;
assign   tb_i_key[532]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[532]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[532]               =   1'b0;
assign   tb_i_rf_static_encrypt[532]          =   1'b1;
assign   tb_i_clear_fault_flags[532]          =   1'b0;
assign   tb_i_rf_static_aad_length[532]       =   64'h0000000000000100;
assign   tb_i_aad[532]                        =   tb_i_aad[531];
assign   tb_i_rf_static_plaintext_length[532] =   64'h0000000000000280;
assign   tb_i_plaintext[532]                  =   tb_i_plaintext[531];
assign   tb_o_valid[532]                      =   1'b0;
assign   tb_o_sop[532]                        =   1'b0;
assign   tb_o_ciphertext[532]                 =   tb_o_ciphertext[531];
assign   tb_o_tag_ready[532]                  =   1'b0;
assign   tb_o_tag[532]                        =   tb_o_tag[531];

// CLK no. 533/1240
// *************************************************
assign   tb_i_valid[533]                      =   1'b1;
assign   tb_i_reset[533]                      =   1'b0;
assign   tb_i_sop[533]                        =   1'b0;
assign   tb_i_key_update[533]                 =   1'b0;
assign   tb_i_key[533]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[533]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[533]               =   1'b0;
assign   tb_i_rf_static_encrypt[533]          =   1'b1;
assign   tb_i_clear_fault_flags[533]          =   1'b0;
assign   tb_i_rf_static_aad_length[533]       =   64'h0000000000000100;
assign   tb_i_aad[533]                        =   256'he6468859a69fb8b20e1a4188090d28946fdfdcf9e193eec9cc906d3f50c2c5ab;
assign   tb_i_rf_static_plaintext_length[533] =   64'h0000000000000280;
assign   tb_i_plaintext[533]                  =   tb_i_plaintext[532];
assign   tb_o_valid[533]                      =   1'b0;
assign   tb_o_sop[533]                        =   1'b0;
assign   tb_o_ciphertext[533]                 =   tb_o_ciphertext[532];
assign   tb_o_tag_ready[533]                  =   1'b0;
assign   tb_o_tag[533]                        =   tb_o_tag[532];

// CLK no. 534/1240
// *************************************************
assign   tb_i_valid[534]                      =   1'b1;
assign   tb_i_reset[534]                      =   1'b0;
assign   tb_i_sop[534]                        =   1'b0;
assign   tb_i_key_update[534]                 =   1'b0;
assign   tb_i_key[534]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[534]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[534]               =   1'b0;
assign   tb_i_rf_static_encrypt[534]          =   1'b1;
assign   tb_i_clear_fault_flags[534]          =   1'b0;
assign   tb_i_rf_static_aad_length[534]       =   64'h0000000000000100;
assign   tb_i_aad[534]                        =   tb_i_aad[533];
assign   tb_i_rf_static_plaintext_length[534] =   64'h0000000000000280;
assign   tb_i_plaintext[534]                  =   256'hec4c20678bbbd6c7445a1421269a7602536150ddafd023c81fb24269a0e9c5aa;
assign   tb_o_valid[534]                      =   1'b0;
assign   tb_o_sop[534]                        =   1'b0;
assign   tb_o_ciphertext[534]                 =   tb_o_ciphertext[533];
assign   tb_o_tag_ready[534]                  =   1'b0;
assign   tb_o_tag[534]                        =   tb_o_tag[533];

// CLK no. 535/1240
// *************************************************
assign   tb_i_valid[535]                      =   1'b1;
assign   tb_i_reset[535]                      =   1'b0;
assign   tb_i_sop[535]                        =   1'b0;
assign   tb_i_key_update[535]                 =   1'b0;
assign   tb_i_key[535]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[535]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[535]               =   1'b0;
assign   tb_i_rf_static_encrypt[535]          =   1'b1;
assign   tb_i_clear_fault_flags[535]          =   1'b0;
assign   tb_i_rf_static_aad_length[535]       =   64'h0000000000000100;
assign   tb_i_aad[535]                        =   tb_i_aad[534];
assign   tb_i_rf_static_plaintext_length[535] =   64'h0000000000000280;
assign   tb_i_plaintext[535]                  =   256'h7d086d01800592ece55419d785ecb881b1f65ffd7d6cf4b73886ad937e8042af;
assign   tb_o_valid[535]                      =   1'b0;
assign   tb_o_sop[535]                        =   1'b0;
assign   tb_o_ciphertext[535]                 =   tb_o_ciphertext[534];
assign   tb_o_tag_ready[535]                  =   1'b0;
assign   tb_o_tag[535]                        =   tb_o_tag[534];

// CLK no. 536/1240
// *************************************************
assign   tb_i_valid[536]                      =   1'b1;
assign   tb_i_reset[536]                      =   1'b0;
assign   tb_i_sop[536]                        =   1'b0;
assign   tb_i_key_update[536]                 =   1'b0;
assign   tb_i_key[536]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[536]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[536]               =   1'b0;
assign   tb_i_rf_static_encrypt[536]          =   1'b1;
assign   tb_i_clear_fault_flags[536]          =   1'b0;
assign   tb_i_rf_static_aad_length[536]       =   64'h0000000000000100;
assign   tb_i_aad[536]                        =   tb_i_aad[535];
assign   tb_i_rf_static_plaintext_length[536] =   64'h0000000000000280;
assign   tb_i_plaintext[536]                  =   256'hae5fc50909dfd6ec490ad9c24141c065;
assign   tb_o_valid[536]                      =   1'b0;
assign   tb_o_sop[536]                        =   1'b0;
assign   tb_o_ciphertext[536]                 =   tb_o_ciphertext[535];
assign   tb_o_tag_ready[536]                  =   1'b0;
assign   tb_o_tag[536]                        =   tb_o_tag[535];

// CLK no. 537/1240
// *************************************************
assign   tb_i_valid[537]                      =   1'b0;
assign   tb_i_reset[537]                      =   1'b0;
assign   tb_i_sop[537]                        =   1'b0;
assign   tb_i_key_update[537]                 =   1'b0;
assign   tb_i_key[537]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[537]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[537]               =   1'b0;
assign   tb_i_rf_static_encrypt[537]          =   1'b1;
assign   tb_i_clear_fault_flags[537]          =   1'b0;
assign   tb_i_rf_static_aad_length[537]       =   64'h0000000000000100;
assign   tb_i_aad[537]                        =   tb_i_aad[536];
assign   tb_i_rf_static_plaintext_length[537] =   64'h0000000000000280;
assign   tb_i_plaintext[537]                  =   tb_i_plaintext[536];
assign   tb_o_valid[537]                      =   1'b0;
assign   tb_o_sop[537]                        =   1'b0;
assign   tb_o_ciphertext[537]                 =   tb_o_ciphertext[536];
assign   tb_o_tag_ready[537]                  =   1'b0;
assign   tb_o_tag[537]                        =   tb_o_tag[536];

// CLK no. 538/1240
// *************************************************
assign   tb_i_valid[538]                      =   1'b0;
assign   tb_i_reset[538]                      =   1'b0;
assign   tb_i_sop[538]                        =   1'b0;
assign   tb_i_key_update[538]                 =   1'b0;
assign   tb_i_key[538]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[538]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[538]               =   1'b0;
assign   tb_i_rf_static_encrypt[538]          =   1'b1;
assign   tb_i_clear_fault_flags[538]          =   1'b0;
assign   tb_i_rf_static_aad_length[538]       =   64'h0000000000000100;
assign   tb_i_aad[538]                        =   tb_i_aad[537];
assign   tb_i_rf_static_plaintext_length[538] =   64'h0000000000000280;
assign   tb_i_plaintext[538]                  =   tb_i_plaintext[537];
assign   tb_o_valid[538]                      =   1'b0;
assign   tb_o_sop[538]                        =   1'b0;
assign   tb_o_ciphertext[538]                 =   tb_o_ciphertext[537];
assign   tb_o_tag_ready[538]                  =   1'b0;
assign   tb_o_tag[538]                        =   tb_o_tag[537];

// CLK no. 539/1240
// *************************************************
assign   tb_i_valid[539]                      =   1'b0;
assign   tb_i_reset[539]                      =   1'b0;
assign   tb_i_sop[539]                        =   1'b0;
assign   tb_i_key_update[539]                 =   1'b0;
assign   tb_i_key[539]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[539]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[539]               =   1'b0;
assign   tb_i_rf_static_encrypt[539]          =   1'b1;
assign   tb_i_clear_fault_flags[539]          =   1'b0;
assign   tb_i_rf_static_aad_length[539]       =   64'h0000000000000100;
assign   tb_i_aad[539]                        =   tb_i_aad[538];
assign   tb_i_rf_static_plaintext_length[539] =   64'h0000000000000280;
assign   tb_i_plaintext[539]                  =   tb_i_plaintext[538];
assign   tb_o_valid[539]                      =   1'b0;
assign   tb_o_sop[539]                        =   1'b0;
assign   tb_o_ciphertext[539]                 =   tb_o_ciphertext[538];
assign   tb_o_tag_ready[539]                  =   1'b0;
assign   tb_o_tag[539]                        =   tb_o_tag[538];

// CLK no. 540/1240
// *************************************************
assign   tb_i_valid[540]                      =   1'b0;
assign   tb_i_reset[540]                      =   1'b0;
assign   tb_i_sop[540]                        =   1'b0;
assign   tb_i_key_update[540]                 =   1'b0;
assign   tb_i_key[540]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[540]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[540]               =   1'b0;
assign   tb_i_rf_static_encrypt[540]          =   1'b1;
assign   tb_i_clear_fault_flags[540]          =   1'b0;
assign   tb_i_rf_static_aad_length[540]       =   64'h0000000000000100;
assign   tb_i_aad[540]                        =   tb_i_aad[539];
assign   tb_i_rf_static_plaintext_length[540] =   64'h0000000000000280;
assign   tb_i_plaintext[540]                  =   tb_i_plaintext[539];
assign   tb_o_valid[540]                      =   1'b0;
assign   tb_o_sop[540]                        =   1'b0;
assign   tb_o_ciphertext[540]                 =   tb_o_ciphertext[539];
assign   tb_o_tag_ready[540]                  =   1'b0;
assign   tb_o_tag[540]                        =   tb_o_tag[539];

// CLK no. 541/1240
// *************************************************
assign   tb_i_valid[541]                      =   1'b0;
assign   tb_i_reset[541]                      =   1'b0;
assign   tb_i_sop[541]                        =   1'b0;
assign   tb_i_key_update[541]                 =   1'b0;
assign   tb_i_key[541]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[541]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[541]               =   1'b0;
assign   tb_i_rf_static_encrypt[541]          =   1'b1;
assign   tb_i_clear_fault_flags[541]          =   1'b0;
assign   tb_i_rf_static_aad_length[541]       =   64'h0000000000000100;
assign   tb_i_aad[541]                        =   tb_i_aad[540];
assign   tb_i_rf_static_plaintext_length[541] =   64'h0000000000000280;
assign   tb_i_plaintext[541]                  =   tb_i_plaintext[540];
assign   tb_o_valid[541]                      =   1'b0;
assign   tb_o_sop[541]                        =   1'b0;
assign   tb_o_ciphertext[541]                 =   tb_o_ciphertext[540];
assign   tb_o_tag_ready[541]                  =   1'b0;
assign   tb_o_tag[541]                        =   tb_o_tag[540];

// CLK no. 542/1240
// *************************************************
assign   tb_i_valid[542]                      =   1'b0;
assign   tb_i_reset[542]                      =   1'b0;
assign   tb_i_sop[542]                        =   1'b0;
assign   tb_i_key_update[542]                 =   1'b0;
assign   tb_i_key[542]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[542]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[542]               =   1'b0;
assign   tb_i_rf_static_encrypt[542]          =   1'b1;
assign   tb_i_clear_fault_flags[542]          =   1'b0;
assign   tb_i_rf_static_aad_length[542]       =   64'h0000000000000100;
assign   tb_i_aad[542]                        =   tb_i_aad[541];
assign   tb_i_rf_static_plaintext_length[542] =   64'h0000000000000280;
assign   tb_i_plaintext[542]                  =   tb_i_plaintext[541];
assign   tb_o_valid[542]                      =   1'b0;
assign   tb_o_sop[542]                        =   1'b0;
assign   tb_o_ciphertext[542]                 =   tb_o_ciphertext[541];
assign   tb_o_tag_ready[542]                  =   1'b0;
assign   tb_o_tag[542]                        =   tb_o_tag[541];

// CLK no. 543/1240
// *************************************************
assign   tb_i_valid[543]                      =   1'b0;
assign   tb_i_reset[543]                      =   1'b0;
assign   tb_i_sop[543]                        =   1'b0;
assign   tb_i_key_update[543]                 =   1'b0;
assign   tb_i_key[543]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[543]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[543]               =   1'b0;
assign   tb_i_rf_static_encrypt[543]          =   1'b1;
assign   tb_i_clear_fault_flags[543]          =   1'b0;
assign   tb_i_rf_static_aad_length[543]       =   64'h0000000000000100;
assign   tb_i_aad[543]                        =   tb_i_aad[542];
assign   tb_i_rf_static_plaintext_length[543] =   64'h0000000000000280;
assign   tb_i_plaintext[543]                  =   tb_i_plaintext[542];
assign   tb_o_valid[543]                      =   1'b0;
assign   tb_o_sop[543]                        =   1'b0;
assign   tb_o_ciphertext[543]                 =   tb_o_ciphertext[542];
assign   tb_o_tag_ready[543]                  =   1'b0;
assign   tb_o_tag[543]                        =   tb_o_tag[542];

// CLK no. 544/1240
// *************************************************
assign   tb_i_valid[544]                      =   1'b0;
assign   tb_i_reset[544]                      =   1'b0;
assign   tb_i_sop[544]                        =   1'b0;
assign   tb_i_key_update[544]                 =   1'b0;
assign   tb_i_key[544]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[544]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[544]               =   1'b0;
assign   tb_i_rf_static_encrypt[544]          =   1'b1;
assign   tb_i_clear_fault_flags[544]          =   1'b0;
assign   tb_i_rf_static_aad_length[544]       =   64'h0000000000000100;
assign   tb_i_aad[544]                        =   tb_i_aad[543];
assign   tb_i_rf_static_plaintext_length[544] =   64'h0000000000000280;
assign   tb_i_plaintext[544]                  =   tb_i_plaintext[543];
assign   tb_o_valid[544]                      =   1'b0;
assign   tb_o_sop[544]                        =   1'b0;
assign   tb_o_ciphertext[544]                 =   tb_o_ciphertext[543];
assign   tb_o_tag_ready[544]                  =   1'b0;
assign   tb_o_tag[544]                        =   tb_o_tag[543];

// CLK no. 545/1240
// *************************************************
assign   tb_i_valid[545]                      =   1'b0;
assign   tb_i_reset[545]                      =   1'b0;
assign   tb_i_sop[545]                        =   1'b0;
assign   tb_i_key_update[545]                 =   1'b0;
assign   tb_i_key[545]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[545]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[545]               =   1'b0;
assign   tb_i_rf_static_encrypt[545]          =   1'b1;
assign   tb_i_clear_fault_flags[545]          =   1'b0;
assign   tb_i_rf_static_aad_length[545]       =   64'h0000000000000100;
assign   tb_i_aad[545]                        =   tb_i_aad[544];
assign   tb_i_rf_static_plaintext_length[545] =   64'h0000000000000280;
assign   tb_i_plaintext[545]                  =   tb_i_plaintext[544];
assign   tb_o_valid[545]                      =   1'b0;
assign   tb_o_sop[545]                        =   1'b0;
assign   tb_o_ciphertext[545]                 =   tb_o_ciphertext[544];
assign   tb_o_tag_ready[545]                  =   1'b0;
assign   tb_o_tag[545]                        =   tb_o_tag[544];

// CLK no. 546/1240
// *************************************************
assign   tb_i_valid[546]                      =   1'b0;
assign   tb_i_reset[546]                      =   1'b0;
assign   tb_i_sop[546]                        =   1'b0;
assign   tb_i_key_update[546]                 =   1'b0;
assign   tb_i_key[546]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[546]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[546]               =   1'b0;
assign   tb_i_rf_static_encrypt[546]          =   1'b1;
assign   tb_i_clear_fault_flags[546]          =   1'b0;
assign   tb_i_rf_static_aad_length[546]       =   64'h0000000000000100;
assign   tb_i_aad[546]                        =   tb_i_aad[545];
assign   tb_i_rf_static_plaintext_length[546] =   64'h0000000000000280;
assign   tb_i_plaintext[546]                  =   tb_i_plaintext[545];
assign   tb_o_valid[546]                      =   1'b0;
assign   tb_o_sop[546]                        =   1'b0;
assign   tb_o_ciphertext[546]                 =   tb_o_ciphertext[545];
assign   tb_o_tag_ready[546]                  =   1'b0;
assign   tb_o_tag[546]                        =   tb_o_tag[545];

// CLK no. 547/1240
// *************************************************
assign   tb_i_valid[547]                      =   1'b0;
assign   tb_i_reset[547]                      =   1'b0;
assign   tb_i_sop[547]                        =   1'b0;
assign   tb_i_key_update[547]                 =   1'b0;
assign   tb_i_key[547]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[547]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[547]               =   1'b0;
assign   tb_i_rf_static_encrypt[547]          =   1'b1;
assign   tb_i_clear_fault_flags[547]          =   1'b0;
assign   tb_i_rf_static_aad_length[547]       =   64'h0000000000000100;
assign   tb_i_aad[547]                        =   tb_i_aad[546];
assign   tb_i_rf_static_plaintext_length[547] =   64'h0000000000000280;
assign   tb_i_plaintext[547]                  =   tb_i_plaintext[546];
assign   tb_o_valid[547]                      =   1'b0;
assign   tb_o_sop[547]                        =   1'b0;
assign   tb_o_ciphertext[547]                 =   tb_o_ciphertext[546];
assign   tb_o_tag_ready[547]                  =   1'b0;
assign   tb_o_tag[547]                        =   tb_o_tag[546];

// CLK no. 548/1240
// *************************************************
assign   tb_i_valid[548]                      =   1'b0;
assign   tb_i_reset[548]                      =   1'b0;
assign   tb_i_sop[548]                        =   1'b0;
assign   tb_i_key_update[548]                 =   1'b0;
assign   tb_i_key[548]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[548]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[548]               =   1'b0;
assign   tb_i_rf_static_encrypt[548]          =   1'b1;
assign   tb_i_clear_fault_flags[548]          =   1'b0;
assign   tb_i_rf_static_aad_length[548]       =   64'h0000000000000100;
assign   tb_i_aad[548]                        =   tb_i_aad[547];
assign   tb_i_rf_static_plaintext_length[548] =   64'h0000000000000280;
assign   tb_i_plaintext[548]                  =   tb_i_plaintext[547];
assign   tb_o_valid[548]                      =   1'b0;
assign   tb_o_sop[548]                        =   1'b0;
assign   tb_o_ciphertext[548]                 =   tb_o_ciphertext[547];
assign   tb_o_tag_ready[548]                  =   1'b0;
assign   tb_o_tag[548]                        =   tb_o_tag[547];

// CLK no. 549/1240
// *************************************************
assign   tb_i_valid[549]                      =   1'b0;
assign   tb_i_reset[549]                      =   1'b0;
assign   tb_i_sop[549]                        =   1'b0;
assign   tb_i_key_update[549]                 =   1'b0;
assign   tb_i_key[549]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[549]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[549]               =   1'b0;
assign   tb_i_rf_static_encrypt[549]          =   1'b1;
assign   tb_i_clear_fault_flags[549]          =   1'b0;
assign   tb_i_rf_static_aad_length[549]       =   64'h0000000000000100;
assign   tb_i_aad[549]                        =   tb_i_aad[548];
assign   tb_i_rf_static_plaintext_length[549] =   64'h0000000000000280;
assign   tb_i_plaintext[549]                  =   tb_i_plaintext[548];
assign   tb_o_valid[549]                      =   1'b0;
assign   tb_o_sop[549]                        =   1'b0;
assign   tb_o_ciphertext[549]                 =   tb_o_ciphertext[548];
assign   tb_o_tag_ready[549]                  =   1'b0;
assign   tb_o_tag[549]                        =   tb_o_tag[548];

// CLK no. 550/1240
// *************************************************
assign   tb_i_valid[550]                      =   1'b0;
assign   tb_i_reset[550]                      =   1'b0;
assign   tb_i_sop[550]                        =   1'b0;
assign   tb_i_key_update[550]                 =   1'b0;
assign   tb_i_key[550]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[550]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[550]               =   1'b0;
assign   tb_i_rf_static_encrypt[550]          =   1'b1;
assign   tb_i_clear_fault_flags[550]          =   1'b0;
assign   tb_i_rf_static_aad_length[550]       =   64'h0000000000000100;
assign   tb_i_aad[550]                        =   tb_i_aad[549];
assign   tb_i_rf_static_plaintext_length[550] =   64'h0000000000000280;
assign   tb_i_plaintext[550]                  =   tb_i_plaintext[549];
assign   tb_o_valid[550]                      =   1'b0;
assign   tb_o_sop[550]                        =   1'b0;
assign   tb_o_ciphertext[550]                 =   tb_o_ciphertext[549];
assign   tb_o_tag_ready[550]                  =   1'b0;
assign   tb_o_tag[550]                        =   tb_o_tag[549];

// CLK no. 551/1240
// *************************************************
assign   tb_i_valid[551]                      =   1'b0;
assign   tb_i_reset[551]                      =   1'b0;
assign   tb_i_sop[551]                        =   1'b0;
assign   tb_i_key_update[551]                 =   1'b0;
assign   tb_i_key[551]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[551]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[551]               =   1'b0;
assign   tb_i_rf_static_encrypt[551]          =   1'b1;
assign   tb_i_clear_fault_flags[551]          =   1'b0;
assign   tb_i_rf_static_aad_length[551]       =   64'h0000000000000100;
assign   tb_i_aad[551]                        =   tb_i_aad[550];
assign   tb_i_rf_static_plaintext_length[551] =   64'h0000000000000280;
assign   tb_i_plaintext[551]                  =   tb_i_plaintext[550];
assign   tb_o_valid[551]                      =   1'b0;
assign   tb_o_sop[551]                        =   1'b0;
assign   tb_o_ciphertext[551]                 =   tb_o_ciphertext[550];
assign   tb_o_tag_ready[551]                  =   1'b0;
assign   tb_o_tag[551]                        =   tb_o_tag[550];

// CLK no. 552/1240
// *************************************************
assign   tb_i_valid[552]                      =   1'b0;
assign   tb_i_reset[552]                      =   1'b0;
assign   tb_i_sop[552]                        =   1'b0;
assign   tb_i_key_update[552]                 =   1'b0;
assign   tb_i_key[552]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[552]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[552]               =   1'b0;
assign   tb_i_rf_static_encrypt[552]          =   1'b1;
assign   tb_i_clear_fault_flags[552]          =   1'b0;
assign   tb_i_rf_static_aad_length[552]       =   64'h0000000000000100;
assign   tb_i_aad[552]                        =   tb_i_aad[551];
assign   tb_i_rf_static_plaintext_length[552] =   64'h0000000000000280;
assign   tb_i_plaintext[552]                  =   tb_i_plaintext[551];
assign   tb_o_valid[552]                      =   1'b0;
assign   tb_o_sop[552]                        =   1'b0;
assign   tb_o_ciphertext[552]                 =   tb_o_ciphertext[551];
assign   tb_o_tag_ready[552]                  =   1'b0;
assign   tb_o_tag[552]                        =   tb_o_tag[551];

// CLK no. 553/1240
// *************************************************
assign   tb_i_valid[553]                      =   1'b0;
assign   tb_i_reset[553]                      =   1'b0;
assign   tb_i_sop[553]                        =   1'b0;
assign   tb_i_key_update[553]                 =   1'b0;
assign   tb_i_key[553]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[553]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[553]               =   1'b0;
assign   tb_i_rf_static_encrypt[553]          =   1'b1;
assign   tb_i_clear_fault_flags[553]          =   1'b0;
assign   tb_i_rf_static_aad_length[553]       =   64'h0000000000000100;
assign   tb_i_aad[553]                        =   tb_i_aad[552];
assign   tb_i_rf_static_plaintext_length[553] =   64'h0000000000000280;
assign   tb_i_plaintext[553]                  =   tb_i_plaintext[552];
assign   tb_o_valid[553]                      =   1'b0;
assign   tb_o_sop[553]                        =   1'b0;
assign   tb_o_ciphertext[553]                 =   tb_o_ciphertext[552];
assign   tb_o_tag_ready[553]                  =   1'b0;
assign   tb_o_tag[553]                        =   tb_o_tag[552];

// CLK no. 554/1240
// *************************************************
assign   tb_i_valid[554]                      =   1'b0;
assign   tb_i_reset[554]                      =   1'b0;
assign   tb_i_sop[554]                        =   1'b0;
assign   tb_i_key_update[554]                 =   1'b0;
assign   tb_i_key[554]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[554]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[554]               =   1'b0;
assign   tb_i_rf_static_encrypt[554]          =   1'b1;
assign   tb_i_clear_fault_flags[554]          =   1'b0;
assign   tb_i_rf_static_aad_length[554]       =   64'h0000000000000100;
assign   tb_i_aad[554]                        =   tb_i_aad[553];
assign   tb_i_rf_static_plaintext_length[554] =   64'h0000000000000280;
assign   tb_i_plaintext[554]                  =   tb_i_plaintext[553];
assign   tb_o_valid[554]                      =   1'b0;
assign   tb_o_sop[554]                        =   1'b0;
assign   tb_o_ciphertext[554]                 =   tb_o_ciphertext[553];
assign   tb_o_tag_ready[554]                  =   1'b0;
assign   tb_o_tag[554]                        =   tb_o_tag[553];

// CLK no. 555/1240
// *************************************************
assign   tb_i_valid[555]                      =   1'b0;
assign   tb_i_reset[555]                      =   1'b0;
assign   tb_i_sop[555]                        =   1'b0;
assign   tb_i_key_update[555]                 =   1'b0;
assign   tb_i_key[555]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[555]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[555]               =   1'b0;
assign   tb_i_rf_static_encrypt[555]          =   1'b1;
assign   tb_i_clear_fault_flags[555]          =   1'b0;
assign   tb_i_rf_static_aad_length[555]       =   64'h0000000000000100;
assign   tb_i_aad[555]                        =   tb_i_aad[554];
assign   tb_i_rf_static_plaintext_length[555] =   64'h0000000000000280;
assign   tb_i_plaintext[555]                  =   tb_i_plaintext[554];
assign   tb_o_valid[555]                      =   1'b0;
assign   tb_o_sop[555]                        =   1'b0;
assign   tb_o_ciphertext[555]                 =   tb_o_ciphertext[554];
assign   tb_o_tag_ready[555]                  =   1'b0;
assign   tb_o_tag[555]                        =   tb_o_tag[554];

// CLK no. 556/1240
// *************************************************
assign   tb_i_valid[556]                      =   1'b0;
assign   tb_i_reset[556]                      =   1'b0;
assign   tb_i_sop[556]                        =   1'b0;
assign   tb_i_key_update[556]                 =   1'b0;
assign   tb_i_key[556]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[556]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[556]               =   1'b0;
assign   tb_i_rf_static_encrypt[556]          =   1'b1;
assign   tb_i_clear_fault_flags[556]          =   1'b0;
assign   tb_i_rf_static_aad_length[556]       =   64'h0000000000000100;
assign   tb_i_aad[556]                        =   tb_i_aad[555];
assign   tb_i_rf_static_plaintext_length[556] =   64'h0000000000000280;
assign   tb_i_plaintext[556]                  =   tb_i_plaintext[555];
assign   tb_o_valid[556]                      =   1'b0;
assign   tb_o_sop[556]                        =   1'b0;
assign   tb_o_ciphertext[556]                 =   tb_o_ciphertext[555];
assign   tb_o_tag_ready[556]                  =   1'b0;
assign   tb_o_tag[556]                        =   tb_o_tag[555];

// CLK no. 557/1240
// *************************************************
assign   tb_i_valid[557]                      =   1'b0;
assign   tb_i_reset[557]                      =   1'b0;
assign   tb_i_sop[557]                        =   1'b0;
assign   tb_i_key_update[557]                 =   1'b0;
assign   tb_i_key[557]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[557]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[557]               =   1'b0;
assign   tb_i_rf_static_encrypt[557]          =   1'b1;
assign   tb_i_clear_fault_flags[557]          =   1'b0;
assign   tb_i_rf_static_aad_length[557]       =   64'h0000000000000100;
assign   tb_i_aad[557]                        =   tb_i_aad[556];
assign   tb_i_rf_static_plaintext_length[557] =   64'h0000000000000280;
assign   tb_i_plaintext[557]                  =   tb_i_plaintext[556];
assign   tb_o_valid[557]                      =   1'b0;
assign   tb_o_sop[557]                        =   1'b0;
assign   tb_o_ciphertext[557]                 =   tb_o_ciphertext[556];
assign   tb_o_tag_ready[557]                  =   1'b0;
assign   tb_o_tag[557]                        =   tb_o_tag[556];

// CLK no. 558/1240
// *************************************************
assign   tb_i_valid[558]                      =   1'b0;
assign   tb_i_reset[558]                      =   1'b0;
assign   tb_i_sop[558]                        =   1'b0;
assign   tb_i_key_update[558]                 =   1'b0;
assign   tb_i_key[558]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[558]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[558]               =   1'b0;
assign   tb_i_rf_static_encrypt[558]          =   1'b1;
assign   tb_i_clear_fault_flags[558]          =   1'b0;
assign   tb_i_rf_static_aad_length[558]       =   64'h0000000000000100;
assign   tb_i_aad[558]                        =   tb_i_aad[557];
assign   tb_i_rf_static_plaintext_length[558] =   64'h0000000000000280;
assign   tb_i_plaintext[558]                  =   tb_i_plaintext[557];
assign   tb_o_valid[558]                      =   1'b0;
assign   tb_o_sop[558]                        =   1'b0;
assign   tb_o_ciphertext[558]                 =   tb_o_ciphertext[557];
assign   tb_o_tag_ready[558]                  =   1'b0;
assign   tb_o_tag[558]                        =   tb_o_tag[557];

// CLK no. 559/1240
// *************************************************
assign   tb_i_valid[559]                      =   1'b0;
assign   tb_i_reset[559]                      =   1'b0;
assign   tb_i_sop[559]                        =   1'b0;
assign   tb_i_key_update[559]                 =   1'b0;
assign   tb_i_key[559]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[559]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[559]               =   1'b0;
assign   tb_i_rf_static_encrypt[559]          =   1'b1;
assign   tb_i_clear_fault_flags[559]          =   1'b0;
assign   tb_i_rf_static_aad_length[559]       =   64'h0000000000000100;
assign   tb_i_aad[559]                        =   tb_i_aad[558];
assign   tb_i_rf_static_plaintext_length[559] =   64'h0000000000000280;
assign   tb_i_plaintext[559]                  =   tb_i_plaintext[558];
assign   tb_o_valid[559]                      =   1'b0;
assign   tb_o_sop[559]                        =   1'b0;
assign   tb_o_ciphertext[559]                 =   tb_o_ciphertext[558];
assign   tb_o_tag_ready[559]                  =   1'b0;
assign   tb_o_tag[559]                        =   tb_o_tag[558];

// CLK no. 560/1240
// *************************************************
assign   tb_i_valid[560]                      =   1'b0;
assign   tb_i_reset[560]                      =   1'b0;
assign   tb_i_sop[560]                        =   1'b0;
assign   tb_i_key_update[560]                 =   1'b0;
assign   tb_i_key[560]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[560]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[560]               =   1'b0;
assign   tb_i_rf_static_encrypt[560]          =   1'b1;
assign   tb_i_clear_fault_flags[560]          =   1'b0;
assign   tb_i_rf_static_aad_length[560]       =   64'h0000000000000100;
assign   tb_i_aad[560]                        =   tb_i_aad[559];
assign   tb_i_rf_static_plaintext_length[560] =   64'h0000000000000280;
assign   tb_i_plaintext[560]                  =   tb_i_plaintext[559];
assign   tb_o_valid[560]                      =   1'b0;
assign   tb_o_sop[560]                        =   1'b0;
assign   tb_o_ciphertext[560]                 =   tb_o_ciphertext[559];
assign   tb_o_tag_ready[560]                  =   1'b0;
assign   tb_o_tag[560]                        =   tb_o_tag[559];

// CLK no. 561/1240
// *************************************************
assign   tb_i_valid[561]                      =   1'b0;
assign   tb_i_reset[561]                      =   1'b0;
assign   tb_i_sop[561]                        =   1'b0;
assign   tb_i_key_update[561]                 =   1'b0;
assign   tb_i_key[561]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[561]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[561]               =   1'b0;
assign   tb_i_rf_static_encrypt[561]          =   1'b1;
assign   tb_i_clear_fault_flags[561]          =   1'b0;
assign   tb_i_rf_static_aad_length[561]       =   64'h0000000000000100;
assign   tb_i_aad[561]                        =   tb_i_aad[560];
assign   tb_i_rf_static_plaintext_length[561] =   64'h0000000000000280;
assign   tb_i_plaintext[561]                  =   tb_i_plaintext[560];
assign   tb_o_valid[561]                      =   1'b0;
assign   tb_o_sop[561]                        =   1'b0;
assign   tb_o_ciphertext[561]                 =   tb_o_ciphertext[560];
assign   tb_o_tag_ready[561]                  =   1'b0;
assign   tb_o_tag[561]                        =   tb_o_tag[560];

// CLK no. 562/1240
// *************************************************
assign   tb_i_valid[562]                      =   1'b0;
assign   tb_i_reset[562]                      =   1'b0;
assign   tb_i_sop[562]                        =   1'b0;
assign   tb_i_key_update[562]                 =   1'b0;
assign   tb_i_key[562]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[562]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[562]               =   1'b0;
assign   tb_i_rf_static_encrypt[562]          =   1'b1;
assign   tb_i_clear_fault_flags[562]          =   1'b0;
assign   tb_i_rf_static_aad_length[562]       =   64'h0000000000000100;
assign   tb_i_aad[562]                        =   tb_i_aad[561];
assign   tb_i_rf_static_plaintext_length[562] =   64'h0000000000000280;
assign   tb_i_plaintext[562]                  =   tb_i_plaintext[561];
assign   tb_o_valid[562]                      =   1'b0;
assign   tb_o_sop[562]                        =   1'b0;
assign   tb_o_ciphertext[562]                 =   tb_o_ciphertext[561];
assign   tb_o_tag_ready[562]                  =   1'b0;
assign   tb_o_tag[562]                        =   tb_o_tag[561];

// CLK no. 563/1240
// *************************************************
assign   tb_i_valid[563]                      =   1'b0;
assign   tb_i_reset[563]                      =   1'b0;
assign   tb_i_sop[563]                        =   1'b0;
assign   tb_i_key_update[563]                 =   1'b0;
assign   tb_i_key[563]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[563]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[563]               =   1'b0;
assign   tb_i_rf_static_encrypt[563]          =   1'b1;
assign   tb_i_clear_fault_flags[563]          =   1'b0;
assign   tb_i_rf_static_aad_length[563]       =   64'h0000000000000100;
assign   tb_i_aad[563]                        =   tb_i_aad[562];
assign   tb_i_rf_static_plaintext_length[563] =   64'h0000000000000280;
assign   tb_i_plaintext[563]                  =   tb_i_plaintext[562];
assign   tb_o_valid[563]                      =   1'b0;
assign   tb_o_sop[563]                        =   1'b0;
assign   tb_o_ciphertext[563]                 =   tb_o_ciphertext[562];
assign   tb_o_tag_ready[563]                  =   1'b0;
assign   tb_o_tag[563]                        =   tb_o_tag[562];

// CLK no. 564/1240
// *************************************************
assign   tb_i_valid[564]                      =   1'b0;
assign   tb_i_reset[564]                      =   1'b0;
assign   tb_i_sop[564]                        =   1'b0;
assign   tb_i_key_update[564]                 =   1'b0;
assign   tb_i_key[564]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[564]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[564]               =   1'b0;
assign   tb_i_rf_static_encrypt[564]          =   1'b1;
assign   tb_i_clear_fault_flags[564]          =   1'b0;
assign   tb_i_rf_static_aad_length[564]       =   64'h0000000000000100;
assign   tb_i_aad[564]                        =   tb_i_aad[563];
assign   tb_i_rf_static_plaintext_length[564] =   64'h0000000000000280;
assign   tb_i_plaintext[564]                  =   tb_i_plaintext[563];
assign   tb_o_valid[564]                      =   1'b0;
assign   tb_o_sop[564]                        =   1'b0;
assign   tb_o_ciphertext[564]                 =   tb_o_ciphertext[563];
assign   tb_o_tag_ready[564]                  =   1'b0;
assign   tb_o_tag[564]                        =   tb_o_tag[563];

// CLK no. 565/1240
// *************************************************
assign   tb_i_valid[565]                      =   1'b0;
assign   tb_i_reset[565]                      =   1'b0;
assign   tb_i_sop[565]                        =   1'b0;
assign   tb_i_key_update[565]                 =   1'b0;
assign   tb_i_key[565]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[565]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[565]               =   1'b0;
assign   tb_i_rf_static_encrypt[565]          =   1'b1;
assign   tb_i_clear_fault_flags[565]          =   1'b0;
assign   tb_i_rf_static_aad_length[565]       =   64'h0000000000000100;
assign   tb_i_aad[565]                        =   tb_i_aad[564];
assign   tb_i_rf_static_plaintext_length[565] =   64'h0000000000000280;
assign   tb_i_plaintext[565]                  =   tb_i_plaintext[564];
assign   tb_o_valid[565]                      =   1'b0;
assign   tb_o_sop[565]                        =   1'b0;
assign   tb_o_ciphertext[565]                 =   tb_o_ciphertext[564];
assign   tb_o_tag_ready[565]                  =   1'b0;
assign   tb_o_tag[565]                        =   tb_o_tag[564];

// CLK no. 566/1240
// *************************************************
assign   tb_i_valid[566]                      =   1'b0;
assign   tb_i_reset[566]                      =   1'b0;
assign   tb_i_sop[566]                        =   1'b0;
assign   tb_i_key_update[566]                 =   1'b0;
assign   tb_i_key[566]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[566]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[566]               =   1'b0;
assign   tb_i_rf_static_encrypt[566]          =   1'b1;
assign   tb_i_clear_fault_flags[566]          =   1'b0;
assign   tb_i_rf_static_aad_length[566]       =   64'h0000000000000100;
assign   tb_i_aad[566]                        =   tb_i_aad[565];
assign   tb_i_rf_static_plaintext_length[566] =   64'h0000000000000280;
assign   tb_i_plaintext[566]                  =   tb_i_plaintext[565];
assign   tb_o_valid[566]                      =   1'b0;
assign   tb_o_sop[566]                        =   1'b0;
assign   tb_o_ciphertext[566]                 =   tb_o_ciphertext[565];
assign   tb_o_tag_ready[566]                  =   1'b0;
assign   tb_o_tag[566]                        =   tb_o_tag[565];

// CLK no. 567/1240
// *************************************************
assign   tb_i_valid[567]                      =   1'b0;
assign   tb_i_reset[567]                      =   1'b0;
assign   tb_i_sop[567]                        =   1'b0;
assign   tb_i_key_update[567]                 =   1'b0;
assign   tb_i_key[567]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[567]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[567]               =   1'b0;
assign   tb_i_rf_static_encrypt[567]          =   1'b1;
assign   tb_i_clear_fault_flags[567]          =   1'b0;
assign   tb_i_rf_static_aad_length[567]       =   64'h0000000000000100;
assign   tb_i_aad[567]                        =   tb_i_aad[566];
assign   tb_i_rf_static_plaintext_length[567] =   64'h0000000000000280;
assign   tb_i_plaintext[567]                  =   tb_i_plaintext[566];
assign   tb_o_valid[567]                      =   1'b0;
assign   tb_o_sop[567]                        =   1'b0;
assign   tb_o_ciphertext[567]                 =   tb_o_ciphertext[566];
assign   tb_o_tag_ready[567]                  =   1'b0;
assign   tb_o_tag[567]                        =   tb_o_tag[566];

// CLK no. 568/1240
// *************************************************
assign   tb_i_valid[568]                      =   1'b0;
assign   tb_i_reset[568]                      =   1'b0;
assign   tb_i_sop[568]                        =   1'b0;
assign   tb_i_key_update[568]                 =   1'b0;
assign   tb_i_key[568]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[568]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[568]               =   1'b0;
assign   tb_i_rf_static_encrypt[568]          =   1'b1;
assign   tb_i_clear_fault_flags[568]          =   1'b0;
assign   tb_i_rf_static_aad_length[568]       =   64'h0000000000000100;
assign   tb_i_aad[568]                        =   tb_i_aad[567];
assign   tb_i_rf_static_plaintext_length[568] =   64'h0000000000000280;
assign   tb_i_plaintext[568]                  =   tb_i_plaintext[567];
assign   tb_o_valid[568]                      =   1'b0;
assign   tb_o_sop[568]                        =   1'b0;
assign   tb_o_ciphertext[568]                 =   tb_o_ciphertext[567];
assign   tb_o_tag_ready[568]                  =   1'b0;
assign   tb_o_tag[568]                        =   tb_o_tag[567];

// CLK no. 569/1240
// *************************************************
assign   tb_i_valid[569]                      =   1'b0;
assign   tb_i_reset[569]                      =   1'b0;
assign   tb_i_sop[569]                        =   1'b0;
assign   tb_i_key_update[569]                 =   1'b0;
assign   tb_i_key[569]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[569]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[569]               =   1'b0;
assign   tb_i_rf_static_encrypt[569]          =   1'b1;
assign   tb_i_clear_fault_flags[569]          =   1'b0;
assign   tb_i_rf_static_aad_length[569]       =   64'h0000000000000100;
assign   tb_i_aad[569]                        =   tb_i_aad[568];
assign   tb_i_rf_static_plaintext_length[569] =   64'h0000000000000280;
assign   tb_i_plaintext[569]                  =   tb_i_plaintext[568];
assign   tb_o_valid[569]                      =   1'b0;
assign   tb_o_sop[569]                        =   1'b0;
assign   tb_o_ciphertext[569]                 =   tb_o_ciphertext[568];
assign   tb_o_tag_ready[569]                  =   1'b0;
assign   tb_o_tag[569]                        =   tb_o_tag[568];

// CLK no. 570/1240
// *************************************************
assign   tb_i_valid[570]                      =   1'b0;
assign   tb_i_reset[570]                      =   1'b0;
assign   tb_i_sop[570]                        =   1'b0;
assign   tb_i_key_update[570]                 =   1'b0;
assign   tb_i_key[570]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[570]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[570]               =   1'b0;
assign   tb_i_rf_static_encrypt[570]          =   1'b1;
assign   tb_i_clear_fault_flags[570]          =   1'b0;
assign   tb_i_rf_static_aad_length[570]       =   64'h0000000000000100;
assign   tb_i_aad[570]                        =   tb_i_aad[569];
assign   tb_i_rf_static_plaintext_length[570] =   64'h0000000000000280;
assign   tb_i_plaintext[570]                  =   tb_i_plaintext[569];
assign   tb_o_valid[570]                      =   1'b0;
assign   tb_o_sop[570]                        =   1'b0;
assign   tb_o_ciphertext[570]                 =   tb_o_ciphertext[569];
assign   tb_o_tag_ready[570]                  =   1'b0;
assign   tb_o_tag[570]                        =   tb_o_tag[569];

// CLK no. 571/1240
// *************************************************
assign   tb_i_valid[571]                      =   1'b0;
assign   tb_i_reset[571]                      =   1'b0;
assign   tb_i_sop[571]                        =   1'b0;
assign   tb_i_key_update[571]                 =   1'b0;
assign   tb_i_key[571]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[571]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[571]               =   1'b0;
assign   tb_i_rf_static_encrypt[571]          =   1'b1;
assign   tb_i_clear_fault_flags[571]          =   1'b0;
assign   tb_i_rf_static_aad_length[571]       =   64'h0000000000000100;
assign   tb_i_aad[571]                        =   tb_i_aad[570];
assign   tb_i_rf_static_plaintext_length[571] =   64'h0000000000000280;
assign   tb_i_plaintext[571]                  =   tb_i_plaintext[570];
assign   tb_o_valid[571]                      =   1'b0;
assign   tb_o_sop[571]                        =   1'b0;
assign   tb_o_ciphertext[571]                 =   tb_o_ciphertext[570];
assign   tb_o_tag_ready[571]                  =   1'b0;
assign   tb_o_tag[571]                        =   tb_o_tag[570];

// CLK no. 572/1240
// *************************************************
assign   tb_i_valid[572]                      =   1'b0;
assign   tb_i_reset[572]                      =   1'b0;
assign   tb_i_sop[572]                        =   1'b0;
assign   tb_i_key_update[572]                 =   1'b0;
assign   tb_i_key[572]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[572]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[572]               =   1'b0;
assign   tb_i_rf_static_encrypt[572]          =   1'b1;
assign   tb_i_clear_fault_flags[572]          =   1'b0;
assign   tb_i_rf_static_aad_length[572]       =   64'h0000000000000100;
assign   tb_i_aad[572]                        =   tb_i_aad[571];
assign   tb_i_rf_static_plaintext_length[572] =   64'h0000000000000280;
assign   tb_i_plaintext[572]                  =   tb_i_plaintext[571];
assign   tb_o_valid[572]                      =   1'b0;
assign   tb_o_sop[572]                        =   1'b0;
assign   tb_o_ciphertext[572]                 =   tb_o_ciphertext[571];
assign   tb_o_tag_ready[572]                  =   1'b0;
assign   tb_o_tag[572]                        =   tb_o_tag[571];

// CLK no. 573/1240
// *************************************************
assign   tb_i_valid[573]                      =   1'b0;
assign   tb_i_reset[573]                      =   1'b0;
assign   tb_i_sop[573]                        =   1'b0;
assign   tb_i_key_update[573]                 =   1'b0;
assign   tb_i_key[573]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[573]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[573]               =   1'b0;
assign   tb_i_rf_static_encrypt[573]          =   1'b1;
assign   tb_i_clear_fault_flags[573]          =   1'b0;
assign   tb_i_rf_static_aad_length[573]       =   64'h0000000000000100;
assign   tb_i_aad[573]                        =   tb_i_aad[572];
assign   tb_i_rf_static_plaintext_length[573] =   64'h0000000000000280;
assign   tb_i_plaintext[573]                  =   tb_i_plaintext[572];
assign   tb_o_valid[573]                      =   1'b0;
assign   tb_o_sop[573]                        =   1'b0;
assign   tb_o_ciphertext[573]                 =   tb_o_ciphertext[572];
assign   tb_o_tag_ready[573]                  =   1'b0;
assign   tb_o_tag[573]                        =   tb_o_tag[572];

// CLK no. 574/1240
// *************************************************
assign   tb_i_valid[574]                      =   1'b0;
assign   tb_i_reset[574]                      =   1'b0;
assign   tb_i_sop[574]                        =   1'b0;
assign   tb_i_key_update[574]                 =   1'b0;
assign   tb_i_key[574]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[574]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[574]               =   1'b0;
assign   tb_i_rf_static_encrypt[574]          =   1'b1;
assign   tb_i_clear_fault_flags[574]          =   1'b0;
assign   tb_i_rf_static_aad_length[574]       =   64'h0000000000000100;
assign   tb_i_aad[574]                        =   tb_i_aad[573];
assign   tb_i_rf_static_plaintext_length[574] =   64'h0000000000000280;
assign   tb_i_plaintext[574]                  =   tb_i_plaintext[573];
assign   tb_o_valid[574]                      =   1'b0;
assign   tb_o_sop[574]                        =   1'b0;
assign   tb_o_ciphertext[574]                 =   tb_o_ciphertext[573];
assign   tb_o_tag_ready[574]                  =   1'b0;
assign   tb_o_tag[574]                        =   tb_o_tag[573];

// CLK no. 575/1240
// *************************************************
assign   tb_i_valid[575]                      =   1'b0;
assign   tb_i_reset[575]                      =   1'b0;
assign   tb_i_sop[575]                        =   1'b0;
assign   tb_i_key_update[575]                 =   1'b0;
assign   tb_i_key[575]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[575]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[575]               =   1'b0;
assign   tb_i_rf_static_encrypt[575]          =   1'b1;
assign   tb_i_clear_fault_flags[575]          =   1'b0;
assign   tb_i_rf_static_aad_length[575]       =   64'h0000000000000100;
assign   tb_i_aad[575]                        =   tb_i_aad[574];
assign   tb_i_rf_static_plaintext_length[575] =   64'h0000000000000280;
assign   tb_i_plaintext[575]                  =   tb_i_plaintext[574];
assign   tb_o_valid[575]                      =   1'b0;
assign   tb_o_sop[575]                        =   1'b0;
assign   tb_o_ciphertext[575]                 =   tb_o_ciphertext[574];
assign   tb_o_tag_ready[575]                  =   1'b0;
assign   tb_o_tag[575]                        =   tb_o_tag[574];

// CLK no. 576/1240
// *************************************************
assign   tb_i_valid[576]                      =   1'b0;
assign   tb_i_reset[576]                      =   1'b0;
assign   tb_i_sop[576]                        =   1'b0;
assign   tb_i_key_update[576]                 =   1'b0;
assign   tb_i_key[576]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[576]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[576]               =   1'b0;
assign   tb_i_rf_static_encrypt[576]          =   1'b1;
assign   tb_i_clear_fault_flags[576]          =   1'b0;
assign   tb_i_rf_static_aad_length[576]       =   64'h0000000000000100;
assign   tb_i_aad[576]                        =   tb_i_aad[575];
assign   tb_i_rf_static_plaintext_length[576] =   64'h0000000000000280;
assign   tb_i_plaintext[576]                  =   tb_i_plaintext[575];
assign   tb_o_valid[576]                      =   1'b0;
assign   tb_o_sop[576]                        =   1'b0;
assign   tb_o_ciphertext[576]                 =   tb_o_ciphertext[575];
assign   tb_o_tag_ready[576]                  =   1'b0;
assign   tb_o_tag[576]                        =   tb_o_tag[575];

// CLK no. 577/1240
// *************************************************
assign   tb_i_valid[577]                      =   1'b0;
assign   tb_i_reset[577]                      =   1'b0;
assign   tb_i_sop[577]                        =   1'b0;
assign   tb_i_key_update[577]                 =   1'b0;
assign   tb_i_key[577]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[577]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[577]               =   1'b0;
assign   tb_i_rf_static_encrypt[577]          =   1'b1;
assign   tb_i_clear_fault_flags[577]          =   1'b0;
assign   tb_i_rf_static_aad_length[577]       =   64'h0000000000000100;
assign   tb_i_aad[577]                        =   tb_i_aad[576];
assign   tb_i_rf_static_plaintext_length[577] =   64'h0000000000000280;
assign   tb_i_plaintext[577]                  =   tb_i_plaintext[576];
assign   tb_o_valid[577]                      =   1'b0;
assign   tb_o_sop[577]                        =   1'b0;
assign   tb_o_ciphertext[577]                 =   tb_o_ciphertext[576];
assign   tb_o_tag_ready[577]                  =   1'b0;
assign   tb_o_tag[577]                        =   tb_o_tag[576];

// CLK no. 578/1240
// *************************************************
assign   tb_i_valid[578]                      =   1'b0;
assign   tb_i_reset[578]                      =   1'b0;
assign   tb_i_sop[578]                        =   1'b0;
assign   tb_i_key_update[578]                 =   1'b0;
assign   tb_i_key[578]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[578]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[578]               =   1'b0;
assign   tb_i_rf_static_encrypt[578]          =   1'b1;
assign   tb_i_clear_fault_flags[578]          =   1'b0;
assign   tb_i_rf_static_aad_length[578]       =   64'h0000000000000100;
assign   tb_i_aad[578]                        =   tb_i_aad[577];
assign   tb_i_rf_static_plaintext_length[578] =   64'h0000000000000280;
assign   tb_i_plaintext[578]                  =   tb_i_plaintext[577];
assign   tb_o_valid[578]                      =   1'b1;
assign   tb_o_sop[578]                        =   1'b1;
assign   tb_o_ciphertext[578]                 =   256'h0ed105e8216ae1d41f8e86a189fe2ddad87da308ce02582a4e947c0f2598a14d;
assign   tb_o_tag_ready[578]                  =   1'b0;
assign   tb_o_tag[578]                        =   tb_o_tag[577];

// CLK no. 579/1240
// *************************************************
assign   tb_i_valid[579]                      =   1'b0;
assign   tb_i_reset[579]                      =   1'b0;
assign   tb_i_sop[579]                        =   1'b0;
assign   tb_i_key_update[579]                 =   1'b0;
assign   tb_i_key[579]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[579]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[579]               =   1'b0;
assign   tb_i_rf_static_encrypt[579]          =   1'b1;
assign   tb_i_clear_fault_flags[579]          =   1'b0;
assign   tb_i_rf_static_aad_length[579]       =   64'h0000000000000100;
assign   tb_i_aad[579]                        =   tb_i_aad[578];
assign   tb_i_rf_static_plaintext_length[579] =   64'h0000000000000280;
assign   tb_i_plaintext[579]                  =   tb_i_plaintext[578];
assign   tb_o_valid[579]                      =   1'b1;
assign   tb_o_sop[579]                        =   1'b0;
assign   tb_o_ciphertext[579]                 =   256'h09949e97b9b20eb1e3fe948c16c37f79217add20b10946d9b0f928a761a47fb2;
assign   tb_o_tag_ready[579]                  =   1'b0;
assign   tb_o_tag[579]                        =   tb_o_tag[578];

// CLK no. 580/1240
// *************************************************
assign   tb_i_valid[580]                      =   1'b0;
assign   tb_i_reset[580]                      =   1'b0;
assign   tb_i_sop[580]                        =   1'b0;
assign   tb_i_key_update[580]                 =   1'b0;
assign   tb_i_key[580]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[580]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[580]               =   1'b0;
assign   tb_i_rf_static_encrypt[580]          =   1'b1;
assign   tb_i_clear_fault_flags[580]          =   1'b0;
assign   tb_i_rf_static_aad_length[580]       =   64'h0000000000000100;
assign   tb_i_aad[580]                        =   tb_i_aad[579];
assign   tb_i_rf_static_plaintext_length[580] =   64'h0000000000000280;
assign   tb_i_plaintext[580]                  =   tb_i_plaintext[579];
assign   tb_o_valid[580]                      =   1'b1;
assign   tb_o_sop[580]                        =   1'b0;
assign   tb_o_ciphertext[580]                 =   256'hcaf0be5fe932aba6019f57dfb7b9208a;
assign   tb_o_tag_ready[580]                  =   1'b0;
assign   tb_o_tag[580]                        =   tb_o_tag[579];

// CLK no. 581/1240
// *************************************************
assign   tb_i_valid[581]                      =   1'b0;
assign   tb_i_reset[581]                      =   1'b0;
assign   tb_i_sop[581]                        =   1'b0;
assign   tb_i_key_update[581]                 =   1'b0;
assign   tb_i_key[581]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[581]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[581]               =   1'b0;
assign   tb_i_rf_static_encrypt[581]          =   1'b1;
assign   tb_i_clear_fault_flags[581]          =   1'b0;
assign   tb_i_rf_static_aad_length[581]       =   64'h0000000000000100;
assign   tb_i_aad[581]                        =   tb_i_aad[580];
assign   tb_i_rf_static_plaintext_length[581] =   64'h0000000000000280;
assign   tb_i_plaintext[581]                  =   tb_i_plaintext[580];
assign   tb_o_valid[581]                      =   1'b0;
assign   tb_o_sop[581]                        =   1'b0;
assign   tb_o_ciphertext[581]                 =   tb_o_ciphertext[580];
assign   tb_o_tag_ready[581]                  =   1'b0;
assign   tb_o_tag[581]                        =   tb_o_tag[580];

// CLK no. 582/1240
// *************************************************
assign   tb_i_valid[582]                      =   1'b0;
assign   tb_i_reset[582]                      =   1'b0;
assign   tb_i_sop[582]                        =   1'b0;
assign   tb_i_key_update[582]                 =   1'b0;
assign   tb_i_key[582]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[582]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[582]               =   1'b0;
assign   tb_i_rf_static_encrypt[582]          =   1'b1;
assign   tb_i_clear_fault_flags[582]          =   1'b0;
assign   tb_i_rf_static_aad_length[582]       =   64'h0000000000000100;
assign   tb_i_aad[582]                        =   tb_i_aad[581];
assign   tb_i_rf_static_plaintext_length[582] =   64'h0000000000000280;
assign   tb_i_plaintext[582]                  =   tb_i_plaintext[581];
assign   tb_o_valid[582]                      =   1'b0;
assign   tb_o_sop[582]                        =   1'b0;
assign   tb_o_ciphertext[582]                 =   tb_o_ciphertext[581];
assign   tb_o_tag_ready[582]                  =   1'b0;
assign   tb_o_tag[582]                        =   tb_o_tag[581];

// CLK no. 583/1240
// *************************************************
assign   tb_i_valid[583]                      =   1'b0;
assign   tb_i_reset[583]                      =   1'b0;
assign   tb_i_sop[583]                        =   1'b0;
assign   tb_i_key_update[583]                 =   1'b0;
assign   tb_i_key[583]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[583]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[583]               =   1'b0;
assign   tb_i_rf_static_encrypt[583]          =   1'b1;
assign   tb_i_clear_fault_flags[583]          =   1'b0;
assign   tb_i_rf_static_aad_length[583]       =   64'h0000000000000100;
assign   tb_i_aad[583]                        =   tb_i_aad[582];
assign   tb_i_rf_static_plaintext_length[583] =   64'h0000000000000280;
assign   tb_i_plaintext[583]                  =   tb_i_plaintext[582];
assign   tb_o_valid[583]                      =   1'b0;
assign   tb_o_sop[583]                        =   1'b0;
assign   tb_o_ciphertext[583]                 =   tb_o_ciphertext[582];
assign   tb_o_tag_ready[583]                  =   1'b0;
assign   tb_o_tag[583]                        =   tb_o_tag[582];

// CLK no. 584/1240
// *************************************************
assign   tb_i_valid[584]                      =   1'b0;
assign   tb_i_reset[584]                      =   1'b0;
assign   tb_i_sop[584]                        =   1'b0;
assign   tb_i_key_update[584]                 =   1'b0;
assign   tb_i_key[584]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[584]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[584]               =   1'b0;
assign   tb_i_rf_static_encrypt[584]          =   1'b1;
assign   tb_i_clear_fault_flags[584]          =   1'b0;
assign   tb_i_rf_static_aad_length[584]       =   64'h0000000000000100;
assign   tb_i_aad[584]                        =   tb_i_aad[583];
assign   tb_i_rf_static_plaintext_length[584] =   64'h0000000000000280;
assign   tb_i_plaintext[584]                  =   tb_i_plaintext[583];
assign   tb_o_valid[584]                      =   1'b0;
assign   tb_o_sop[584]                        =   1'b0;
assign   tb_o_ciphertext[584]                 =   tb_o_ciphertext[583];
assign   tb_o_tag_ready[584]                  =   1'b0;
assign   tb_o_tag[584]                        =   tb_o_tag[583];

// CLK no. 585/1240
// *************************************************
assign   tb_i_valid[585]                      =   1'b0;
assign   tb_i_reset[585]                      =   1'b0;
assign   tb_i_sop[585]                        =   1'b0;
assign   tb_i_key_update[585]                 =   1'b0;
assign   tb_i_key[585]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[585]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[585]               =   1'b0;
assign   tb_i_rf_static_encrypt[585]          =   1'b1;
assign   tb_i_clear_fault_flags[585]          =   1'b0;
assign   tb_i_rf_static_aad_length[585]       =   64'h0000000000000100;
assign   tb_i_aad[585]                        =   tb_i_aad[584];
assign   tb_i_rf_static_plaintext_length[585] =   64'h0000000000000280;
assign   tb_i_plaintext[585]                  =   tb_i_plaintext[584];
assign   tb_o_valid[585]                      =   1'b0;
assign   tb_o_sop[585]                        =   1'b0;
assign   tb_o_ciphertext[585]                 =   tb_o_ciphertext[584];
assign   tb_o_tag_ready[585]                  =   1'b0;
assign   tb_o_tag[585]                        =   tb_o_tag[584];

// CLK no. 586/1240
// *************************************************
assign   tb_i_valid[586]                      =   1'b0;
assign   tb_i_reset[586]                      =   1'b0;
assign   tb_i_sop[586]                        =   1'b0;
assign   tb_i_key_update[586]                 =   1'b0;
assign   tb_i_key[586]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[586]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[586]               =   1'b0;
assign   tb_i_rf_static_encrypt[586]          =   1'b1;
assign   tb_i_clear_fault_flags[586]          =   1'b0;
assign   tb_i_rf_static_aad_length[586]       =   64'h0000000000000100;
assign   tb_i_aad[586]                        =   tb_i_aad[585];
assign   tb_i_rf_static_plaintext_length[586] =   64'h0000000000000280;
assign   tb_i_plaintext[586]                  =   tb_i_plaintext[585];
assign   tb_o_valid[586]                      =   1'b0;
assign   tb_o_sop[586]                        =   1'b0;
assign   tb_o_ciphertext[586]                 =   tb_o_ciphertext[585];
assign   tb_o_tag_ready[586]                  =   1'b0;
assign   tb_o_tag[586]                        =   tb_o_tag[585];

// CLK no. 587/1240
// *************************************************
assign   tb_i_valid[587]                      =   1'b0;
assign   tb_i_reset[587]                      =   1'b0;
assign   tb_i_sop[587]                        =   1'b0;
assign   tb_i_key_update[587]                 =   1'b0;
assign   tb_i_key[587]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[587]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[587]               =   1'b0;
assign   tb_i_rf_static_encrypt[587]          =   1'b1;
assign   tb_i_clear_fault_flags[587]          =   1'b0;
assign   tb_i_rf_static_aad_length[587]       =   64'h0000000000000100;
assign   tb_i_aad[587]                        =   tb_i_aad[586];
assign   tb_i_rf_static_plaintext_length[587] =   64'h0000000000000280;
assign   tb_i_plaintext[587]                  =   tb_i_plaintext[586];
assign   tb_o_valid[587]                      =   1'b0;
assign   tb_o_sop[587]                        =   1'b0;
assign   tb_o_ciphertext[587]                 =   tb_o_ciphertext[586];
assign   tb_o_tag_ready[587]                  =   1'b0;
assign   tb_o_tag[587]                        =   tb_o_tag[586];

// CLK no. 588/1240
// *************************************************
assign   tb_i_valid[588]                      =   1'b0;
assign   tb_i_reset[588]                      =   1'b0;
assign   tb_i_sop[588]                        =   1'b0;
assign   tb_i_key_update[588]                 =   1'b0;
assign   tb_i_key[588]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[588]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[588]               =   1'b0;
assign   tb_i_rf_static_encrypt[588]          =   1'b1;
assign   tb_i_clear_fault_flags[588]          =   1'b0;
assign   tb_i_rf_static_aad_length[588]       =   64'h0000000000000100;
assign   tb_i_aad[588]                        =   tb_i_aad[587];
assign   tb_i_rf_static_plaintext_length[588] =   64'h0000000000000280;
assign   tb_i_plaintext[588]                  =   tb_i_plaintext[587];
assign   tb_o_valid[588]                      =   1'b0;
assign   tb_o_sop[588]                        =   1'b0;
assign   tb_o_ciphertext[588]                 =   tb_o_ciphertext[587];
assign   tb_o_tag_ready[588]                  =   1'b1;
assign   tb_o_tag[588]                        =   128'hea7982afa83ac6894172051e90b31d04;

// CLK no. 589/1240
// *************************************************
assign   tb_i_valid[589]                      =   1'b0;
assign   tb_i_reset[589]                      =   1'b0;
assign   tb_i_sop[589]                        =   1'b0;
assign   tb_i_key_update[589]                 =   1'b0;
assign   tb_i_key[589]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[589]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[589]               =   1'b0;
assign   tb_i_rf_static_encrypt[589]          =   1'b1;
assign   tb_i_clear_fault_flags[589]          =   1'b0;
assign   tb_i_rf_static_aad_length[589]       =   64'h0000000000000100;
assign   tb_i_aad[589]                        =   tb_i_aad[588];
assign   tb_i_rf_static_plaintext_length[589] =   64'h0000000000000280;
assign   tb_i_plaintext[589]                  =   tb_i_plaintext[588];
assign   tb_o_valid[589]                      =   1'b0;
assign   tb_o_sop[589]                        =   1'b0;
assign   tb_o_ciphertext[589]                 =   tb_o_ciphertext[588];
assign   tb_o_tag_ready[589]                  =   1'b0;
assign   tb_o_tag[589]                        =   tb_o_tag[588];

// CLK no. 590/1240
// *************************************************
assign   tb_i_valid[590]                      =   1'b0;
assign   tb_i_reset[590]                      =   1'b0;
assign   tb_i_sop[590]                        =   1'b0;
assign   tb_i_key_update[590]                 =   1'b0;
assign   tb_i_key[590]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[590]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[590]               =   1'b0;
assign   tb_i_rf_static_encrypt[590]          =   1'b1;
assign   tb_i_clear_fault_flags[590]          =   1'b0;
assign   tb_i_rf_static_aad_length[590]       =   64'h0000000000000100;
assign   tb_i_aad[590]                        =   tb_i_aad[589];
assign   tb_i_rf_static_plaintext_length[590] =   64'h0000000000000280;
assign   tb_i_plaintext[590]                  =   tb_i_plaintext[589];
assign   tb_o_valid[590]                      =   1'b0;
assign   tb_o_sop[590]                        =   1'b0;
assign   tb_o_ciphertext[590]                 =   tb_o_ciphertext[589];
assign   tb_o_tag_ready[590]                  =   1'b0;
assign   tb_o_tag[590]                        =   tb_o_tag[589];

// CLK no. 591/1240
// *************************************************
assign   tb_i_valid[591]                      =   1'b0;
assign   tb_i_reset[591]                      =   1'b0;
assign   tb_i_sop[591]                        =   1'b1;
assign   tb_i_key_update[591]                 =   1'b0;
assign   tb_i_key[591]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[591]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[591]               =   1'b0;
assign   tb_i_rf_static_encrypt[591]          =   1'b1;
assign   tb_i_clear_fault_flags[591]          =   1'b0;
assign   tb_i_rf_static_aad_length[591]       =   64'h0000000000000100;
assign   tb_i_aad[591]                        =   tb_i_aad[590];
assign   tb_i_rf_static_plaintext_length[591] =   64'h0000000000000280;
assign   tb_i_plaintext[591]                  =   tb_i_plaintext[590];
assign   tb_o_valid[591]                      =   1'b0;
assign   tb_o_sop[591]                        =   1'b0;
assign   tb_o_ciphertext[591]                 =   tb_o_ciphertext[590];
assign   tb_o_tag_ready[591]                  =   1'b0;
assign   tb_o_tag[591]                        =   tb_o_tag[590];

// CLK no. 592/1240
// *************************************************
assign   tb_i_valid[592]                      =   1'b1;
assign   tb_i_reset[592]                      =   1'b0;
assign   tb_i_sop[592]                        =   1'b0;
assign   tb_i_key_update[592]                 =   1'b0;
assign   tb_i_key[592]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[592]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[592]               =   1'b0;
assign   tb_i_rf_static_encrypt[592]          =   1'b1;
assign   tb_i_clear_fault_flags[592]          =   1'b0;
assign   tb_i_rf_static_aad_length[592]       =   64'h0000000000000100;
assign   tb_i_aad[592]                        =   256'hff924ec64dac4646fe027142d8cd68bb87daf302b10e6ea29fd2a309d6df7e92;
assign   tb_i_rf_static_plaintext_length[592] =   64'h0000000000000280;
assign   tb_i_plaintext[592]                  =   tb_i_plaintext[591];
assign   tb_o_valid[592]                      =   1'b0;
assign   tb_o_sop[592]                        =   1'b0;
assign   tb_o_ciphertext[592]                 =   tb_o_ciphertext[591];
assign   tb_o_tag_ready[592]                  =   1'b0;
assign   tb_o_tag[592]                        =   tb_o_tag[591];

// CLK no. 593/1240
// *************************************************
assign   tb_i_valid[593]                      =   1'b1;
assign   tb_i_reset[593]                      =   1'b0;
assign   tb_i_sop[593]                        =   1'b0;
assign   tb_i_key_update[593]                 =   1'b0;
assign   tb_i_key[593]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[593]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[593]               =   1'b0;
assign   tb_i_rf_static_encrypt[593]          =   1'b1;
assign   tb_i_clear_fault_flags[593]          =   1'b0;
assign   tb_i_rf_static_aad_length[593]       =   64'h0000000000000100;
assign   tb_i_aad[593]                        =   tb_i_aad[592];
assign   tb_i_rf_static_plaintext_length[593] =   64'h0000000000000280;
assign   tb_i_plaintext[593]                  =   256'h5198810a8afe0d35b372db1a7831ba3d0255a1a51776c1108c6e615899028270;
assign   tb_o_valid[593]                      =   1'b0;
assign   tb_o_sop[593]                        =   1'b0;
assign   tb_o_ciphertext[593]                 =   tb_o_ciphertext[592];
assign   tb_o_tag_ready[593]                  =   1'b0;
assign   tb_o_tag[593]                        =   tb_o_tag[592];

// CLK no. 594/1240
// *************************************************
assign   tb_i_valid[594]                      =   1'b1;
assign   tb_i_reset[594]                      =   1'b0;
assign   tb_i_sop[594]                        =   1'b0;
assign   tb_i_key_update[594]                 =   1'b0;
assign   tb_i_key[594]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[594]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[594]               =   1'b0;
assign   tb_i_rf_static_encrypt[594]          =   1'b1;
assign   tb_i_clear_fault_flags[594]          =   1'b0;
assign   tb_i_rf_static_aad_length[594]       =   64'h0000000000000100;
assign   tb_i_aad[594]                        =   tb_i_aad[593];
assign   tb_i_rf_static_plaintext_length[594] =   64'h0000000000000280;
assign   tb_i_plaintext[594]                  =   256'hc353871a1b7a1b8a4f47b73f74ff3e48bebe13d7fad7f076a47f61fc398f5da2;
assign   tb_o_valid[594]                      =   1'b0;
assign   tb_o_sop[594]                        =   1'b0;
assign   tb_o_ciphertext[594]                 =   tb_o_ciphertext[593];
assign   tb_o_tag_ready[594]                  =   1'b0;
assign   tb_o_tag[594]                        =   tb_o_tag[593];

// CLK no. 595/1240
// *************************************************
assign   tb_i_valid[595]                      =   1'b1;
assign   tb_i_reset[595]                      =   1'b0;
assign   tb_i_sop[595]                        =   1'b0;
assign   tb_i_key_update[595]                 =   1'b0;
assign   tb_i_key[595]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[595]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[595]               =   1'b0;
assign   tb_i_rf_static_encrypt[595]          =   1'b1;
assign   tb_i_clear_fault_flags[595]          =   1'b0;
assign   tb_i_rf_static_aad_length[595]       =   64'h0000000000000100;
assign   tb_i_aad[595]                        =   tb_i_aad[594];
assign   tb_i_rf_static_plaintext_length[595] =   64'h0000000000000280;
assign   tb_i_plaintext[595]                  =   256'hec91e807f1f7df837224f71835aef519;
assign   tb_o_valid[595]                      =   1'b0;
assign   tb_o_sop[595]                        =   1'b0;
assign   tb_o_ciphertext[595]                 =   tb_o_ciphertext[594];
assign   tb_o_tag_ready[595]                  =   1'b0;
assign   tb_o_tag[595]                        =   tb_o_tag[594];

// CLK no. 596/1240
// *************************************************
assign   tb_i_valid[596]                      =   1'b0;
assign   tb_i_reset[596]                      =   1'b0;
assign   tb_i_sop[596]                        =   1'b0;
assign   tb_i_key_update[596]                 =   1'b0;
assign   tb_i_key[596]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[596]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[596]               =   1'b0;
assign   tb_i_rf_static_encrypt[596]          =   1'b1;
assign   tb_i_clear_fault_flags[596]          =   1'b0;
assign   tb_i_rf_static_aad_length[596]       =   64'h0000000000000100;
assign   tb_i_aad[596]                        =   tb_i_aad[595];
assign   tb_i_rf_static_plaintext_length[596] =   64'h0000000000000280;
assign   tb_i_plaintext[596]                  =   tb_i_plaintext[595];
assign   tb_o_valid[596]                      =   1'b0;
assign   tb_o_sop[596]                        =   1'b0;
assign   tb_o_ciphertext[596]                 =   tb_o_ciphertext[595];
assign   tb_o_tag_ready[596]                  =   1'b0;
assign   tb_o_tag[596]                        =   tb_o_tag[595];

// CLK no. 597/1240
// *************************************************
assign   tb_i_valid[597]                      =   1'b0;
assign   tb_i_reset[597]                      =   1'b0;
assign   tb_i_sop[597]                        =   1'b0;
assign   tb_i_key_update[597]                 =   1'b0;
assign   tb_i_key[597]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[597]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[597]               =   1'b0;
assign   tb_i_rf_static_encrypt[597]          =   1'b1;
assign   tb_i_clear_fault_flags[597]          =   1'b0;
assign   tb_i_rf_static_aad_length[597]       =   64'h0000000000000100;
assign   tb_i_aad[597]                        =   tb_i_aad[596];
assign   tb_i_rf_static_plaintext_length[597] =   64'h0000000000000280;
assign   tb_i_plaintext[597]                  =   tb_i_plaintext[596];
assign   tb_o_valid[597]                      =   1'b0;
assign   tb_o_sop[597]                        =   1'b0;
assign   tb_o_ciphertext[597]                 =   tb_o_ciphertext[596];
assign   tb_o_tag_ready[597]                  =   1'b0;
assign   tb_o_tag[597]                        =   tb_o_tag[596];

// CLK no. 598/1240
// *************************************************
assign   tb_i_valid[598]                      =   1'b0;
assign   tb_i_reset[598]                      =   1'b0;
assign   tb_i_sop[598]                        =   1'b0;
assign   tb_i_key_update[598]                 =   1'b0;
assign   tb_i_key[598]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[598]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[598]               =   1'b0;
assign   tb_i_rf_static_encrypt[598]          =   1'b1;
assign   tb_i_clear_fault_flags[598]          =   1'b0;
assign   tb_i_rf_static_aad_length[598]       =   64'h0000000000000100;
assign   tb_i_aad[598]                        =   tb_i_aad[597];
assign   tb_i_rf_static_plaintext_length[598] =   64'h0000000000000280;
assign   tb_i_plaintext[598]                  =   tb_i_plaintext[597];
assign   tb_o_valid[598]                      =   1'b0;
assign   tb_o_sop[598]                        =   1'b0;
assign   tb_o_ciphertext[598]                 =   tb_o_ciphertext[597];
assign   tb_o_tag_ready[598]                  =   1'b0;
assign   tb_o_tag[598]                        =   tb_o_tag[597];

// CLK no. 599/1240
// *************************************************
assign   tb_i_valid[599]                      =   1'b0;
assign   tb_i_reset[599]                      =   1'b0;
assign   tb_i_sop[599]                        =   1'b0;
assign   tb_i_key_update[599]                 =   1'b0;
assign   tb_i_key[599]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[599]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[599]               =   1'b0;
assign   tb_i_rf_static_encrypt[599]          =   1'b1;
assign   tb_i_clear_fault_flags[599]          =   1'b0;
assign   tb_i_rf_static_aad_length[599]       =   64'h0000000000000100;
assign   tb_i_aad[599]                        =   tb_i_aad[598];
assign   tb_i_rf_static_plaintext_length[599] =   64'h0000000000000280;
assign   tb_i_plaintext[599]                  =   tb_i_plaintext[598];
assign   tb_o_valid[599]                      =   1'b0;
assign   tb_o_sop[599]                        =   1'b0;
assign   tb_o_ciphertext[599]                 =   tb_o_ciphertext[598];
assign   tb_o_tag_ready[599]                  =   1'b0;
assign   tb_o_tag[599]                        =   tb_o_tag[598];

// CLK no. 600/1240
// *************************************************
assign   tb_i_valid[600]                      =   1'b0;
assign   tb_i_reset[600]                      =   1'b0;
assign   tb_i_sop[600]                        =   1'b0;
assign   tb_i_key_update[600]                 =   1'b0;
assign   tb_i_key[600]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[600]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[600]               =   1'b0;
assign   tb_i_rf_static_encrypt[600]          =   1'b1;
assign   tb_i_clear_fault_flags[600]          =   1'b0;
assign   tb_i_rf_static_aad_length[600]       =   64'h0000000000000100;
assign   tb_i_aad[600]                        =   tb_i_aad[599];
assign   tb_i_rf_static_plaintext_length[600] =   64'h0000000000000280;
assign   tb_i_plaintext[600]                  =   tb_i_plaintext[599];
assign   tb_o_valid[600]                      =   1'b0;
assign   tb_o_sop[600]                        =   1'b0;
assign   tb_o_ciphertext[600]                 =   tb_o_ciphertext[599];
assign   tb_o_tag_ready[600]                  =   1'b0;
assign   tb_o_tag[600]                        =   tb_o_tag[599];

// CLK no. 601/1240
// *************************************************
assign   tb_i_valid[601]                      =   1'b0;
assign   tb_i_reset[601]                      =   1'b0;
assign   tb_i_sop[601]                        =   1'b0;
assign   tb_i_key_update[601]                 =   1'b0;
assign   tb_i_key[601]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[601]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[601]               =   1'b0;
assign   tb_i_rf_static_encrypt[601]          =   1'b1;
assign   tb_i_clear_fault_flags[601]          =   1'b0;
assign   tb_i_rf_static_aad_length[601]       =   64'h0000000000000100;
assign   tb_i_aad[601]                        =   tb_i_aad[600];
assign   tb_i_rf_static_plaintext_length[601] =   64'h0000000000000280;
assign   tb_i_plaintext[601]                  =   tb_i_plaintext[600];
assign   tb_o_valid[601]                      =   1'b0;
assign   tb_o_sop[601]                        =   1'b0;
assign   tb_o_ciphertext[601]                 =   tb_o_ciphertext[600];
assign   tb_o_tag_ready[601]                  =   1'b0;
assign   tb_o_tag[601]                        =   tb_o_tag[600];

// CLK no. 602/1240
// *************************************************
assign   tb_i_valid[602]                      =   1'b0;
assign   tb_i_reset[602]                      =   1'b0;
assign   tb_i_sop[602]                        =   1'b0;
assign   tb_i_key_update[602]                 =   1'b0;
assign   tb_i_key[602]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[602]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[602]               =   1'b0;
assign   tb_i_rf_static_encrypt[602]          =   1'b1;
assign   tb_i_clear_fault_flags[602]          =   1'b0;
assign   tb_i_rf_static_aad_length[602]       =   64'h0000000000000100;
assign   tb_i_aad[602]                        =   tb_i_aad[601];
assign   tb_i_rf_static_plaintext_length[602] =   64'h0000000000000280;
assign   tb_i_plaintext[602]                  =   tb_i_plaintext[601];
assign   tb_o_valid[602]                      =   1'b0;
assign   tb_o_sop[602]                        =   1'b0;
assign   tb_o_ciphertext[602]                 =   tb_o_ciphertext[601];
assign   tb_o_tag_ready[602]                  =   1'b0;
assign   tb_o_tag[602]                        =   tb_o_tag[601];

// CLK no. 603/1240
// *************************************************
assign   tb_i_valid[603]                      =   1'b0;
assign   tb_i_reset[603]                      =   1'b0;
assign   tb_i_sop[603]                        =   1'b0;
assign   tb_i_key_update[603]                 =   1'b0;
assign   tb_i_key[603]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[603]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[603]               =   1'b0;
assign   tb_i_rf_static_encrypt[603]          =   1'b1;
assign   tb_i_clear_fault_flags[603]          =   1'b0;
assign   tb_i_rf_static_aad_length[603]       =   64'h0000000000000100;
assign   tb_i_aad[603]                        =   tb_i_aad[602];
assign   tb_i_rf_static_plaintext_length[603] =   64'h0000000000000280;
assign   tb_i_plaintext[603]                  =   tb_i_plaintext[602];
assign   tb_o_valid[603]                      =   1'b0;
assign   tb_o_sop[603]                        =   1'b0;
assign   tb_o_ciphertext[603]                 =   tb_o_ciphertext[602];
assign   tb_o_tag_ready[603]                  =   1'b0;
assign   tb_o_tag[603]                        =   tb_o_tag[602];

// CLK no. 604/1240
// *************************************************
assign   tb_i_valid[604]                      =   1'b0;
assign   tb_i_reset[604]                      =   1'b0;
assign   tb_i_sop[604]                        =   1'b0;
assign   tb_i_key_update[604]                 =   1'b0;
assign   tb_i_key[604]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[604]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[604]               =   1'b0;
assign   tb_i_rf_static_encrypt[604]          =   1'b1;
assign   tb_i_clear_fault_flags[604]          =   1'b0;
assign   tb_i_rf_static_aad_length[604]       =   64'h0000000000000100;
assign   tb_i_aad[604]                        =   tb_i_aad[603];
assign   tb_i_rf_static_plaintext_length[604] =   64'h0000000000000280;
assign   tb_i_plaintext[604]                  =   tb_i_plaintext[603];
assign   tb_o_valid[604]                      =   1'b0;
assign   tb_o_sop[604]                        =   1'b0;
assign   tb_o_ciphertext[604]                 =   tb_o_ciphertext[603];
assign   tb_o_tag_ready[604]                  =   1'b0;
assign   tb_o_tag[604]                        =   tb_o_tag[603];

// CLK no. 605/1240
// *************************************************
assign   tb_i_valid[605]                      =   1'b0;
assign   tb_i_reset[605]                      =   1'b0;
assign   tb_i_sop[605]                        =   1'b0;
assign   tb_i_key_update[605]                 =   1'b0;
assign   tb_i_key[605]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[605]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[605]               =   1'b0;
assign   tb_i_rf_static_encrypt[605]          =   1'b1;
assign   tb_i_clear_fault_flags[605]          =   1'b0;
assign   tb_i_rf_static_aad_length[605]       =   64'h0000000000000100;
assign   tb_i_aad[605]                        =   tb_i_aad[604];
assign   tb_i_rf_static_plaintext_length[605] =   64'h0000000000000280;
assign   tb_i_plaintext[605]                  =   tb_i_plaintext[604];
assign   tb_o_valid[605]                      =   1'b0;
assign   tb_o_sop[605]                        =   1'b0;
assign   tb_o_ciphertext[605]                 =   tb_o_ciphertext[604];
assign   tb_o_tag_ready[605]                  =   1'b0;
assign   tb_o_tag[605]                        =   tb_o_tag[604];

// CLK no. 606/1240
// *************************************************
assign   tb_i_valid[606]                      =   1'b0;
assign   tb_i_reset[606]                      =   1'b0;
assign   tb_i_sop[606]                        =   1'b0;
assign   tb_i_key_update[606]                 =   1'b0;
assign   tb_i_key[606]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[606]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[606]               =   1'b0;
assign   tb_i_rf_static_encrypt[606]          =   1'b1;
assign   tb_i_clear_fault_flags[606]          =   1'b0;
assign   tb_i_rf_static_aad_length[606]       =   64'h0000000000000100;
assign   tb_i_aad[606]                        =   tb_i_aad[605];
assign   tb_i_rf_static_plaintext_length[606] =   64'h0000000000000280;
assign   tb_i_plaintext[606]                  =   tb_i_plaintext[605];
assign   tb_o_valid[606]                      =   1'b0;
assign   tb_o_sop[606]                        =   1'b0;
assign   tb_o_ciphertext[606]                 =   tb_o_ciphertext[605];
assign   tb_o_tag_ready[606]                  =   1'b0;
assign   tb_o_tag[606]                        =   tb_o_tag[605];

// CLK no. 607/1240
// *************************************************
assign   tb_i_valid[607]                      =   1'b0;
assign   tb_i_reset[607]                      =   1'b0;
assign   tb_i_sop[607]                        =   1'b0;
assign   tb_i_key_update[607]                 =   1'b0;
assign   tb_i_key[607]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[607]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[607]               =   1'b0;
assign   tb_i_rf_static_encrypt[607]          =   1'b1;
assign   tb_i_clear_fault_flags[607]          =   1'b0;
assign   tb_i_rf_static_aad_length[607]       =   64'h0000000000000100;
assign   tb_i_aad[607]                        =   tb_i_aad[606];
assign   tb_i_rf_static_plaintext_length[607] =   64'h0000000000000280;
assign   tb_i_plaintext[607]                  =   tb_i_plaintext[606];
assign   tb_o_valid[607]                      =   1'b0;
assign   tb_o_sop[607]                        =   1'b0;
assign   tb_o_ciphertext[607]                 =   tb_o_ciphertext[606];
assign   tb_o_tag_ready[607]                  =   1'b0;
assign   tb_o_tag[607]                        =   tb_o_tag[606];

// CLK no. 608/1240
// *************************************************
assign   tb_i_valid[608]                      =   1'b0;
assign   tb_i_reset[608]                      =   1'b0;
assign   tb_i_sop[608]                        =   1'b0;
assign   tb_i_key_update[608]                 =   1'b0;
assign   tb_i_key[608]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[608]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[608]               =   1'b0;
assign   tb_i_rf_static_encrypt[608]          =   1'b1;
assign   tb_i_clear_fault_flags[608]          =   1'b0;
assign   tb_i_rf_static_aad_length[608]       =   64'h0000000000000100;
assign   tb_i_aad[608]                        =   tb_i_aad[607];
assign   tb_i_rf_static_plaintext_length[608] =   64'h0000000000000280;
assign   tb_i_plaintext[608]                  =   tb_i_plaintext[607];
assign   tb_o_valid[608]                      =   1'b0;
assign   tb_o_sop[608]                        =   1'b0;
assign   tb_o_ciphertext[608]                 =   tb_o_ciphertext[607];
assign   tb_o_tag_ready[608]                  =   1'b0;
assign   tb_o_tag[608]                        =   tb_o_tag[607];

// CLK no. 609/1240
// *************************************************
assign   tb_i_valid[609]                      =   1'b0;
assign   tb_i_reset[609]                      =   1'b0;
assign   tb_i_sop[609]                        =   1'b0;
assign   tb_i_key_update[609]                 =   1'b0;
assign   tb_i_key[609]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[609]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[609]               =   1'b0;
assign   tb_i_rf_static_encrypt[609]          =   1'b1;
assign   tb_i_clear_fault_flags[609]          =   1'b0;
assign   tb_i_rf_static_aad_length[609]       =   64'h0000000000000100;
assign   tb_i_aad[609]                        =   tb_i_aad[608];
assign   tb_i_rf_static_plaintext_length[609] =   64'h0000000000000280;
assign   tb_i_plaintext[609]                  =   tb_i_plaintext[608];
assign   tb_o_valid[609]                      =   1'b0;
assign   tb_o_sop[609]                        =   1'b0;
assign   tb_o_ciphertext[609]                 =   tb_o_ciphertext[608];
assign   tb_o_tag_ready[609]                  =   1'b0;
assign   tb_o_tag[609]                        =   tb_o_tag[608];

// CLK no. 610/1240
// *************************************************
assign   tb_i_valid[610]                      =   1'b0;
assign   tb_i_reset[610]                      =   1'b0;
assign   tb_i_sop[610]                        =   1'b0;
assign   tb_i_key_update[610]                 =   1'b0;
assign   tb_i_key[610]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[610]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[610]               =   1'b0;
assign   tb_i_rf_static_encrypt[610]          =   1'b1;
assign   tb_i_clear_fault_flags[610]          =   1'b0;
assign   tb_i_rf_static_aad_length[610]       =   64'h0000000000000100;
assign   tb_i_aad[610]                        =   tb_i_aad[609];
assign   tb_i_rf_static_plaintext_length[610] =   64'h0000000000000280;
assign   tb_i_plaintext[610]                  =   tb_i_plaintext[609];
assign   tb_o_valid[610]                      =   1'b0;
assign   tb_o_sop[610]                        =   1'b0;
assign   tb_o_ciphertext[610]                 =   tb_o_ciphertext[609];
assign   tb_o_tag_ready[610]                  =   1'b0;
assign   tb_o_tag[610]                        =   tb_o_tag[609];

// CLK no. 611/1240
// *************************************************
assign   tb_i_valid[611]                      =   1'b0;
assign   tb_i_reset[611]                      =   1'b0;
assign   tb_i_sop[611]                        =   1'b0;
assign   tb_i_key_update[611]                 =   1'b0;
assign   tb_i_key[611]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[611]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[611]               =   1'b0;
assign   tb_i_rf_static_encrypt[611]          =   1'b1;
assign   tb_i_clear_fault_flags[611]          =   1'b0;
assign   tb_i_rf_static_aad_length[611]       =   64'h0000000000000100;
assign   tb_i_aad[611]                        =   tb_i_aad[610];
assign   tb_i_rf_static_plaintext_length[611] =   64'h0000000000000280;
assign   tb_i_plaintext[611]                  =   tb_i_plaintext[610];
assign   tb_o_valid[611]                      =   1'b0;
assign   tb_o_sop[611]                        =   1'b0;
assign   tb_o_ciphertext[611]                 =   tb_o_ciphertext[610];
assign   tb_o_tag_ready[611]                  =   1'b0;
assign   tb_o_tag[611]                        =   tb_o_tag[610];

// CLK no. 612/1240
// *************************************************
assign   tb_i_valid[612]                      =   1'b0;
assign   tb_i_reset[612]                      =   1'b0;
assign   tb_i_sop[612]                        =   1'b0;
assign   tb_i_key_update[612]                 =   1'b0;
assign   tb_i_key[612]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[612]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[612]               =   1'b0;
assign   tb_i_rf_static_encrypt[612]          =   1'b1;
assign   tb_i_clear_fault_flags[612]          =   1'b0;
assign   tb_i_rf_static_aad_length[612]       =   64'h0000000000000100;
assign   tb_i_aad[612]                        =   tb_i_aad[611];
assign   tb_i_rf_static_plaintext_length[612] =   64'h0000000000000280;
assign   tb_i_plaintext[612]                  =   tb_i_plaintext[611];
assign   tb_o_valid[612]                      =   1'b0;
assign   tb_o_sop[612]                        =   1'b0;
assign   tb_o_ciphertext[612]                 =   tb_o_ciphertext[611];
assign   tb_o_tag_ready[612]                  =   1'b0;
assign   tb_o_tag[612]                        =   tb_o_tag[611];

// CLK no. 613/1240
// *************************************************
assign   tb_i_valid[613]                      =   1'b0;
assign   tb_i_reset[613]                      =   1'b0;
assign   tb_i_sop[613]                        =   1'b0;
assign   tb_i_key_update[613]                 =   1'b0;
assign   tb_i_key[613]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[613]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[613]               =   1'b0;
assign   tb_i_rf_static_encrypt[613]          =   1'b1;
assign   tb_i_clear_fault_flags[613]          =   1'b0;
assign   tb_i_rf_static_aad_length[613]       =   64'h0000000000000100;
assign   tb_i_aad[613]                        =   tb_i_aad[612];
assign   tb_i_rf_static_plaintext_length[613] =   64'h0000000000000280;
assign   tb_i_plaintext[613]                  =   tb_i_plaintext[612];
assign   tb_o_valid[613]                      =   1'b0;
assign   tb_o_sop[613]                        =   1'b0;
assign   tb_o_ciphertext[613]                 =   tb_o_ciphertext[612];
assign   tb_o_tag_ready[613]                  =   1'b0;
assign   tb_o_tag[613]                        =   tb_o_tag[612];

// CLK no. 614/1240
// *************************************************
assign   tb_i_valid[614]                      =   1'b0;
assign   tb_i_reset[614]                      =   1'b0;
assign   tb_i_sop[614]                        =   1'b0;
assign   tb_i_key_update[614]                 =   1'b0;
assign   tb_i_key[614]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[614]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[614]               =   1'b0;
assign   tb_i_rf_static_encrypt[614]          =   1'b1;
assign   tb_i_clear_fault_flags[614]          =   1'b0;
assign   tb_i_rf_static_aad_length[614]       =   64'h0000000000000100;
assign   tb_i_aad[614]                        =   tb_i_aad[613];
assign   tb_i_rf_static_plaintext_length[614] =   64'h0000000000000280;
assign   tb_i_plaintext[614]                  =   tb_i_plaintext[613];
assign   tb_o_valid[614]                      =   1'b0;
assign   tb_o_sop[614]                        =   1'b0;
assign   tb_o_ciphertext[614]                 =   tb_o_ciphertext[613];
assign   tb_o_tag_ready[614]                  =   1'b0;
assign   tb_o_tag[614]                        =   tb_o_tag[613];

// CLK no. 615/1240
// *************************************************
assign   tb_i_valid[615]                      =   1'b0;
assign   tb_i_reset[615]                      =   1'b0;
assign   tb_i_sop[615]                        =   1'b0;
assign   tb_i_key_update[615]                 =   1'b0;
assign   tb_i_key[615]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[615]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[615]               =   1'b0;
assign   tb_i_rf_static_encrypt[615]          =   1'b1;
assign   tb_i_clear_fault_flags[615]          =   1'b0;
assign   tb_i_rf_static_aad_length[615]       =   64'h0000000000000100;
assign   tb_i_aad[615]                        =   tb_i_aad[614];
assign   tb_i_rf_static_plaintext_length[615] =   64'h0000000000000280;
assign   tb_i_plaintext[615]                  =   tb_i_plaintext[614];
assign   tb_o_valid[615]                      =   1'b0;
assign   tb_o_sop[615]                        =   1'b0;
assign   tb_o_ciphertext[615]                 =   tb_o_ciphertext[614];
assign   tb_o_tag_ready[615]                  =   1'b0;
assign   tb_o_tag[615]                        =   tb_o_tag[614];

// CLK no. 616/1240
// *************************************************
assign   tb_i_valid[616]                      =   1'b0;
assign   tb_i_reset[616]                      =   1'b0;
assign   tb_i_sop[616]                        =   1'b0;
assign   tb_i_key_update[616]                 =   1'b0;
assign   tb_i_key[616]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[616]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[616]               =   1'b0;
assign   tb_i_rf_static_encrypt[616]          =   1'b1;
assign   tb_i_clear_fault_flags[616]          =   1'b0;
assign   tb_i_rf_static_aad_length[616]       =   64'h0000000000000100;
assign   tb_i_aad[616]                        =   tb_i_aad[615];
assign   tb_i_rf_static_plaintext_length[616] =   64'h0000000000000280;
assign   tb_i_plaintext[616]                  =   tb_i_plaintext[615];
assign   tb_o_valid[616]                      =   1'b0;
assign   tb_o_sop[616]                        =   1'b0;
assign   tb_o_ciphertext[616]                 =   tb_o_ciphertext[615];
assign   tb_o_tag_ready[616]                  =   1'b0;
assign   tb_o_tag[616]                        =   tb_o_tag[615];

// CLK no. 617/1240
// *************************************************
assign   tb_i_valid[617]                      =   1'b0;
assign   tb_i_reset[617]                      =   1'b0;
assign   tb_i_sop[617]                        =   1'b0;
assign   tb_i_key_update[617]                 =   1'b0;
assign   tb_i_key[617]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[617]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[617]               =   1'b0;
assign   tb_i_rf_static_encrypt[617]          =   1'b1;
assign   tb_i_clear_fault_flags[617]          =   1'b0;
assign   tb_i_rf_static_aad_length[617]       =   64'h0000000000000100;
assign   tb_i_aad[617]                        =   tb_i_aad[616];
assign   tb_i_rf_static_plaintext_length[617] =   64'h0000000000000280;
assign   tb_i_plaintext[617]                  =   tb_i_plaintext[616];
assign   tb_o_valid[617]                      =   1'b0;
assign   tb_o_sop[617]                        =   1'b0;
assign   tb_o_ciphertext[617]                 =   tb_o_ciphertext[616];
assign   tb_o_tag_ready[617]                  =   1'b0;
assign   tb_o_tag[617]                        =   tb_o_tag[616];

// CLK no. 618/1240
// *************************************************
assign   tb_i_valid[618]                      =   1'b0;
assign   tb_i_reset[618]                      =   1'b0;
assign   tb_i_sop[618]                        =   1'b0;
assign   tb_i_key_update[618]                 =   1'b0;
assign   tb_i_key[618]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[618]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[618]               =   1'b0;
assign   tb_i_rf_static_encrypt[618]          =   1'b1;
assign   tb_i_clear_fault_flags[618]          =   1'b0;
assign   tb_i_rf_static_aad_length[618]       =   64'h0000000000000100;
assign   tb_i_aad[618]                        =   tb_i_aad[617];
assign   tb_i_rf_static_plaintext_length[618] =   64'h0000000000000280;
assign   tb_i_plaintext[618]                  =   tb_i_plaintext[617];
assign   tb_o_valid[618]                      =   1'b0;
assign   tb_o_sop[618]                        =   1'b0;
assign   tb_o_ciphertext[618]                 =   tb_o_ciphertext[617];
assign   tb_o_tag_ready[618]                  =   1'b0;
assign   tb_o_tag[618]                        =   tb_o_tag[617];

// CLK no. 619/1240
// *************************************************
assign   tb_i_valid[619]                      =   1'b0;
assign   tb_i_reset[619]                      =   1'b0;
assign   tb_i_sop[619]                        =   1'b0;
assign   tb_i_key_update[619]                 =   1'b0;
assign   tb_i_key[619]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[619]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[619]               =   1'b0;
assign   tb_i_rf_static_encrypt[619]          =   1'b1;
assign   tb_i_clear_fault_flags[619]          =   1'b0;
assign   tb_i_rf_static_aad_length[619]       =   64'h0000000000000100;
assign   tb_i_aad[619]                        =   tb_i_aad[618];
assign   tb_i_rf_static_plaintext_length[619] =   64'h0000000000000280;
assign   tb_i_plaintext[619]                  =   tb_i_plaintext[618];
assign   tb_o_valid[619]                      =   1'b0;
assign   tb_o_sop[619]                        =   1'b0;
assign   tb_o_ciphertext[619]                 =   tb_o_ciphertext[618];
assign   tb_o_tag_ready[619]                  =   1'b0;
assign   tb_o_tag[619]                        =   tb_o_tag[618];

// CLK no. 620/1240
// *************************************************
assign   tb_i_valid[620]                      =   1'b0;
assign   tb_i_reset[620]                      =   1'b0;
assign   tb_i_sop[620]                        =   1'b0;
assign   tb_i_key_update[620]                 =   1'b0;
assign   tb_i_key[620]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[620]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[620]               =   1'b0;
assign   tb_i_rf_static_encrypt[620]          =   1'b1;
assign   tb_i_clear_fault_flags[620]          =   1'b0;
assign   tb_i_rf_static_aad_length[620]       =   64'h0000000000000100;
assign   tb_i_aad[620]                        =   tb_i_aad[619];
assign   tb_i_rf_static_plaintext_length[620] =   64'h0000000000000280;
assign   tb_i_plaintext[620]                  =   tb_i_plaintext[619];
assign   tb_o_valid[620]                      =   1'b0;
assign   tb_o_sop[620]                        =   1'b0;
assign   tb_o_ciphertext[620]                 =   tb_o_ciphertext[619];
assign   tb_o_tag_ready[620]                  =   1'b0;
assign   tb_o_tag[620]                        =   tb_o_tag[619];

// CLK no. 621/1240
// *************************************************
assign   tb_i_valid[621]                      =   1'b0;
assign   tb_i_reset[621]                      =   1'b0;
assign   tb_i_sop[621]                        =   1'b0;
assign   tb_i_key_update[621]                 =   1'b0;
assign   tb_i_key[621]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[621]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[621]               =   1'b0;
assign   tb_i_rf_static_encrypt[621]          =   1'b1;
assign   tb_i_clear_fault_flags[621]          =   1'b0;
assign   tb_i_rf_static_aad_length[621]       =   64'h0000000000000100;
assign   tb_i_aad[621]                        =   tb_i_aad[620];
assign   tb_i_rf_static_plaintext_length[621] =   64'h0000000000000280;
assign   tb_i_plaintext[621]                  =   tb_i_plaintext[620];
assign   tb_o_valid[621]                      =   1'b0;
assign   tb_o_sop[621]                        =   1'b0;
assign   tb_o_ciphertext[621]                 =   tb_o_ciphertext[620];
assign   tb_o_tag_ready[621]                  =   1'b0;
assign   tb_o_tag[621]                        =   tb_o_tag[620];

// CLK no. 622/1240
// *************************************************
assign   tb_i_valid[622]                      =   1'b0;
assign   tb_i_reset[622]                      =   1'b0;
assign   tb_i_sop[622]                        =   1'b0;
assign   tb_i_key_update[622]                 =   1'b0;
assign   tb_i_key[622]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[622]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[622]               =   1'b0;
assign   tb_i_rf_static_encrypt[622]          =   1'b1;
assign   tb_i_clear_fault_flags[622]          =   1'b0;
assign   tb_i_rf_static_aad_length[622]       =   64'h0000000000000100;
assign   tb_i_aad[622]                        =   tb_i_aad[621];
assign   tb_i_rf_static_plaintext_length[622] =   64'h0000000000000280;
assign   tb_i_plaintext[622]                  =   tb_i_plaintext[621];
assign   tb_o_valid[622]                      =   1'b0;
assign   tb_o_sop[622]                        =   1'b0;
assign   tb_o_ciphertext[622]                 =   tb_o_ciphertext[621];
assign   tb_o_tag_ready[622]                  =   1'b0;
assign   tb_o_tag[622]                        =   tb_o_tag[621];

// CLK no. 623/1240
// *************************************************
assign   tb_i_valid[623]                      =   1'b0;
assign   tb_i_reset[623]                      =   1'b0;
assign   tb_i_sop[623]                        =   1'b0;
assign   tb_i_key_update[623]                 =   1'b0;
assign   tb_i_key[623]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[623]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[623]               =   1'b0;
assign   tb_i_rf_static_encrypt[623]          =   1'b1;
assign   tb_i_clear_fault_flags[623]          =   1'b0;
assign   tb_i_rf_static_aad_length[623]       =   64'h0000000000000100;
assign   tb_i_aad[623]                        =   tb_i_aad[622];
assign   tb_i_rf_static_plaintext_length[623] =   64'h0000000000000280;
assign   tb_i_plaintext[623]                  =   tb_i_plaintext[622];
assign   tb_o_valid[623]                      =   1'b0;
assign   tb_o_sop[623]                        =   1'b0;
assign   tb_o_ciphertext[623]                 =   tb_o_ciphertext[622];
assign   tb_o_tag_ready[623]                  =   1'b0;
assign   tb_o_tag[623]                        =   tb_o_tag[622];

// CLK no. 624/1240
// *************************************************
assign   tb_i_valid[624]                      =   1'b0;
assign   tb_i_reset[624]                      =   1'b0;
assign   tb_i_sop[624]                        =   1'b0;
assign   tb_i_key_update[624]                 =   1'b0;
assign   tb_i_key[624]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[624]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[624]               =   1'b0;
assign   tb_i_rf_static_encrypt[624]          =   1'b1;
assign   tb_i_clear_fault_flags[624]          =   1'b0;
assign   tb_i_rf_static_aad_length[624]       =   64'h0000000000000100;
assign   tb_i_aad[624]                        =   tb_i_aad[623];
assign   tb_i_rf_static_plaintext_length[624] =   64'h0000000000000280;
assign   tb_i_plaintext[624]                  =   tb_i_plaintext[623];
assign   tb_o_valid[624]                      =   1'b0;
assign   tb_o_sop[624]                        =   1'b0;
assign   tb_o_ciphertext[624]                 =   tb_o_ciphertext[623];
assign   tb_o_tag_ready[624]                  =   1'b0;
assign   tb_o_tag[624]                        =   tb_o_tag[623];

// CLK no. 625/1240
// *************************************************
assign   tb_i_valid[625]                      =   1'b0;
assign   tb_i_reset[625]                      =   1'b0;
assign   tb_i_sop[625]                        =   1'b0;
assign   tb_i_key_update[625]                 =   1'b0;
assign   tb_i_key[625]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[625]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[625]               =   1'b0;
assign   tb_i_rf_static_encrypt[625]          =   1'b1;
assign   tb_i_clear_fault_flags[625]          =   1'b0;
assign   tb_i_rf_static_aad_length[625]       =   64'h0000000000000100;
assign   tb_i_aad[625]                        =   tb_i_aad[624];
assign   tb_i_rf_static_plaintext_length[625] =   64'h0000000000000280;
assign   tb_i_plaintext[625]                  =   tb_i_plaintext[624];
assign   tb_o_valid[625]                      =   1'b0;
assign   tb_o_sop[625]                        =   1'b0;
assign   tb_o_ciphertext[625]                 =   tb_o_ciphertext[624];
assign   tb_o_tag_ready[625]                  =   1'b0;
assign   tb_o_tag[625]                        =   tb_o_tag[624];

// CLK no. 626/1240
// *************************************************
assign   tb_i_valid[626]                      =   1'b0;
assign   tb_i_reset[626]                      =   1'b0;
assign   tb_i_sop[626]                        =   1'b0;
assign   tb_i_key_update[626]                 =   1'b0;
assign   tb_i_key[626]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[626]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[626]               =   1'b0;
assign   tb_i_rf_static_encrypt[626]          =   1'b1;
assign   tb_i_clear_fault_flags[626]          =   1'b0;
assign   tb_i_rf_static_aad_length[626]       =   64'h0000000000000100;
assign   tb_i_aad[626]                        =   tb_i_aad[625];
assign   tb_i_rf_static_plaintext_length[626] =   64'h0000000000000280;
assign   tb_i_plaintext[626]                  =   tb_i_plaintext[625];
assign   tb_o_valid[626]                      =   1'b0;
assign   tb_o_sop[626]                        =   1'b0;
assign   tb_o_ciphertext[626]                 =   tb_o_ciphertext[625];
assign   tb_o_tag_ready[626]                  =   1'b0;
assign   tb_o_tag[626]                        =   tb_o_tag[625];

// CLK no. 627/1240
// *************************************************
assign   tb_i_valid[627]                      =   1'b0;
assign   tb_i_reset[627]                      =   1'b0;
assign   tb_i_sop[627]                        =   1'b0;
assign   tb_i_key_update[627]                 =   1'b0;
assign   tb_i_key[627]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[627]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[627]               =   1'b0;
assign   tb_i_rf_static_encrypt[627]          =   1'b1;
assign   tb_i_clear_fault_flags[627]          =   1'b0;
assign   tb_i_rf_static_aad_length[627]       =   64'h0000000000000100;
assign   tb_i_aad[627]                        =   tb_i_aad[626];
assign   tb_i_rf_static_plaintext_length[627] =   64'h0000000000000280;
assign   tb_i_plaintext[627]                  =   tb_i_plaintext[626];
assign   tb_o_valid[627]                      =   1'b0;
assign   tb_o_sop[627]                        =   1'b0;
assign   tb_o_ciphertext[627]                 =   tb_o_ciphertext[626];
assign   tb_o_tag_ready[627]                  =   1'b0;
assign   tb_o_tag[627]                        =   tb_o_tag[626];

// CLK no. 628/1240
// *************************************************
assign   tb_i_valid[628]                      =   1'b0;
assign   tb_i_reset[628]                      =   1'b0;
assign   tb_i_sop[628]                        =   1'b0;
assign   tb_i_key_update[628]                 =   1'b0;
assign   tb_i_key[628]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[628]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[628]               =   1'b0;
assign   tb_i_rf_static_encrypt[628]          =   1'b1;
assign   tb_i_clear_fault_flags[628]          =   1'b0;
assign   tb_i_rf_static_aad_length[628]       =   64'h0000000000000100;
assign   tb_i_aad[628]                        =   tb_i_aad[627];
assign   tb_i_rf_static_plaintext_length[628] =   64'h0000000000000280;
assign   tb_i_plaintext[628]                  =   tb_i_plaintext[627];
assign   tb_o_valid[628]                      =   1'b0;
assign   tb_o_sop[628]                        =   1'b0;
assign   tb_o_ciphertext[628]                 =   tb_o_ciphertext[627];
assign   tb_o_tag_ready[628]                  =   1'b0;
assign   tb_o_tag[628]                        =   tb_o_tag[627];

// CLK no. 629/1240
// *************************************************
assign   tb_i_valid[629]                      =   1'b0;
assign   tb_i_reset[629]                      =   1'b0;
assign   tb_i_sop[629]                        =   1'b0;
assign   tb_i_key_update[629]                 =   1'b0;
assign   tb_i_key[629]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[629]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[629]               =   1'b0;
assign   tb_i_rf_static_encrypt[629]          =   1'b1;
assign   tb_i_clear_fault_flags[629]          =   1'b0;
assign   tb_i_rf_static_aad_length[629]       =   64'h0000000000000100;
assign   tb_i_aad[629]                        =   tb_i_aad[628];
assign   tb_i_rf_static_plaintext_length[629] =   64'h0000000000000280;
assign   tb_i_plaintext[629]                  =   tb_i_plaintext[628];
assign   tb_o_valid[629]                      =   1'b0;
assign   tb_o_sop[629]                        =   1'b0;
assign   tb_o_ciphertext[629]                 =   tb_o_ciphertext[628];
assign   tb_o_tag_ready[629]                  =   1'b0;
assign   tb_o_tag[629]                        =   tb_o_tag[628];

// CLK no. 630/1240
// *************************************************
assign   tb_i_valid[630]                      =   1'b0;
assign   tb_i_reset[630]                      =   1'b0;
assign   tb_i_sop[630]                        =   1'b0;
assign   tb_i_key_update[630]                 =   1'b0;
assign   tb_i_key[630]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[630]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[630]               =   1'b0;
assign   tb_i_rf_static_encrypt[630]          =   1'b1;
assign   tb_i_clear_fault_flags[630]          =   1'b0;
assign   tb_i_rf_static_aad_length[630]       =   64'h0000000000000100;
assign   tb_i_aad[630]                        =   tb_i_aad[629];
assign   tb_i_rf_static_plaintext_length[630] =   64'h0000000000000280;
assign   tb_i_plaintext[630]                  =   tb_i_plaintext[629];
assign   tb_o_valid[630]                      =   1'b0;
assign   tb_o_sop[630]                        =   1'b0;
assign   tb_o_ciphertext[630]                 =   tb_o_ciphertext[629];
assign   tb_o_tag_ready[630]                  =   1'b0;
assign   tb_o_tag[630]                        =   tb_o_tag[629];

// CLK no. 631/1240
// *************************************************
assign   tb_i_valid[631]                      =   1'b0;
assign   tb_i_reset[631]                      =   1'b0;
assign   tb_i_sop[631]                        =   1'b0;
assign   tb_i_key_update[631]                 =   1'b0;
assign   tb_i_key[631]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[631]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[631]               =   1'b0;
assign   tb_i_rf_static_encrypt[631]          =   1'b1;
assign   tb_i_clear_fault_flags[631]          =   1'b0;
assign   tb_i_rf_static_aad_length[631]       =   64'h0000000000000100;
assign   tb_i_aad[631]                        =   tb_i_aad[630];
assign   tb_i_rf_static_plaintext_length[631] =   64'h0000000000000280;
assign   tb_i_plaintext[631]                  =   tb_i_plaintext[630];
assign   tb_o_valid[631]                      =   1'b0;
assign   tb_o_sop[631]                        =   1'b0;
assign   tb_o_ciphertext[631]                 =   tb_o_ciphertext[630];
assign   tb_o_tag_ready[631]                  =   1'b0;
assign   tb_o_tag[631]                        =   tb_o_tag[630];

// CLK no. 632/1240
// *************************************************
assign   tb_i_valid[632]                      =   1'b0;
assign   tb_i_reset[632]                      =   1'b0;
assign   tb_i_sop[632]                        =   1'b0;
assign   tb_i_key_update[632]                 =   1'b0;
assign   tb_i_key[632]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[632]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[632]               =   1'b0;
assign   tb_i_rf_static_encrypt[632]          =   1'b1;
assign   tb_i_clear_fault_flags[632]          =   1'b0;
assign   tb_i_rf_static_aad_length[632]       =   64'h0000000000000100;
assign   tb_i_aad[632]                        =   tb_i_aad[631];
assign   tb_i_rf_static_plaintext_length[632] =   64'h0000000000000280;
assign   tb_i_plaintext[632]                  =   tb_i_plaintext[631];
assign   tb_o_valid[632]                      =   1'b0;
assign   tb_o_sop[632]                        =   1'b0;
assign   tb_o_ciphertext[632]                 =   tb_o_ciphertext[631];
assign   tb_o_tag_ready[632]                  =   1'b0;
assign   tb_o_tag[632]                        =   tb_o_tag[631];

// CLK no. 633/1240
// *************************************************
assign   tb_i_valid[633]                      =   1'b0;
assign   tb_i_reset[633]                      =   1'b0;
assign   tb_i_sop[633]                        =   1'b0;
assign   tb_i_key_update[633]                 =   1'b0;
assign   tb_i_key[633]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[633]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[633]               =   1'b0;
assign   tb_i_rf_static_encrypt[633]          =   1'b1;
assign   tb_i_clear_fault_flags[633]          =   1'b0;
assign   tb_i_rf_static_aad_length[633]       =   64'h0000000000000100;
assign   tb_i_aad[633]                        =   tb_i_aad[632];
assign   tb_i_rf_static_plaintext_length[633] =   64'h0000000000000280;
assign   tb_i_plaintext[633]                  =   tb_i_plaintext[632];
assign   tb_o_valid[633]                      =   1'b0;
assign   tb_o_sop[633]                        =   1'b0;
assign   tb_o_ciphertext[633]                 =   tb_o_ciphertext[632];
assign   tb_o_tag_ready[633]                  =   1'b0;
assign   tb_o_tag[633]                        =   tb_o_tag[632];

// CLK no. 634/1240
// *************************************************
assign   tb_i_valid[634]                      =   1'b0;
assign   tb_i_reset[634]                      =   1'b0;
assign   tb_i_sop[634]                        =   1'b0;
assign   tb_i_key_update[634]                 =   1'b0;
assign   tb_i_key[634]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[634]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[634]               =   1'b0;
assign   tb_i_rf_static_encrypt[634]          =   1'b1;
assign   tb_i_clear_fault_flags[634]          =   1'b0;
assign   tb_i_rf_static_aad_length[634]       =   64'h0000000000000100;
assign   tb_i_aad[634]                        =   tb_i_aad[633];
assign   tb_i_rf_static_plaintext_length[634] =   64'h0000000000000280;
assign   tb_i_plaintext[634]                  =   tb_i_plaintext[633];
assign   tb_o_valid[634]                      =   1'b0;
assign   tb_o_sop[634]                        =   1'b0;
assign   tb_o_ciphertext[634]                 =   tb_o_ciphertext[633];
assign   tb_o_tag_ready[634]                  =   1'b0;
assign   tb_o_tag[634]                        =   tb_o_tag[633];

// CLK no. 635/1240
// *************************************************
assign   tb_i_valid[635]                      =   1'b0;
assign   tb_i_reset[635]                      =   1'b0;
assign   tb_i_sop[635]                        =   1'b0;
assign   tb_i_key_update[635]                 =   1'b0;
assign   tb_i_key[635]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[635]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[635]               =   1'b0;
assign   tb_i_rf_static_encrypt[635]          =   1'b1;
assign   tb_i_clear_fault_flags[635]          =   1'b0;
assign   tb_i_rf_static_aad_length[635]       =   64'h0000000000000100;
assign   tb_i_aad[635]                        =   tb_i_aad[634];
assign   tb_i_rf_static_plaintext_length[635] =   64'h0000000000000280;
assign   tb_i_plaintext[635]                  =   tb_i_plaintext[634];
assign   tb_o_valid[635]                      =   1'b0;
assign   tb_o_sop[635]                        =   1'b0;
assign   tb_o_ciphertext[635]                 =   tb_o_ciphertext[634];
assign   tb_o_tag_ready[635]                  =   1'b0;
assign   tb_o_tag[635]                        =   tb_o_tag[634];

// CLK no. 636/1240
// *************************************************
assign   tb_i_valid[636]                      =   1'b0;
assign   tb_i_reset[636]                      =   1'b0;
assign   tb_i_sop[636]                        =   1'b0;
assign   tb_i_key_update[636]                 =   1'b0;
assign   tb_i_key[636]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[636]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[636]               =   1'b0;
assign   tb_i_rf_static_encrypt[636]          =   1'b1;
assign   tb_i_clear_fault_flags[636]          =   1'b0;
assign   tb_i_rf_static_aad_length[636]       =   64'h0000000000000100;
assign   tb_i_aad[636]                        =   tb_i_aad[635];
assign   tb_i_rf_static_plaintext_length[636] =   64'h0000000000000280;
assign   tb_i_plaintext[636]                  =   tb_i_plaintext[635];
assign   tb_o_valid[636]                      =   1'b0;
assign   tb_o_sop[636]                        =   1'b0;
assign   tb_o_ciphertext[636]                 =   tb_o_ciphertext[635];
assign   tb_o_tag_ready[636]                  =   1'b0;
assign   tb_o_tag[636]                        =   tb_o_tag[635];

// CLK no. 637/1240
// *************************************************
assign   tb_i_valid[637]                      =   1'b0;
assign   tb_i_reset[637]                      =   1'b0;
assign   tb_i_sop[637]                        =   1'b0;
assign   tb_i_key_update[637]                 =   1'b0;
assign   tb_i_key[637]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[637]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[637]               =   1'b0;
assign   tb_i_rf_static_encrypt[637]          =   1'b1;
assign   tb_i_clear_fault_flags[637]          =   1'b0;
assign   tb_i_rf_static_aad_length[637]       =   64'h0000000000000100;
assign   tb_i_aad[637]                        =   tb_i_aad[636];
assign   tb_i_rf_static_plaintext_length[637] =   64'h0000000000000280;
assign   tb_i_plaintext[637]                  =   tb_i_plaintext[636];
assign   tb_o_valid[637]                      =   1'b1;
assign   tb_o_sop[637]                        =   1'b1;
assign   tb_o_ciphertext[637]                 =   256'hb305a485202f3a26e8a6499ad755e1e58949527076a4baf2dd485f3e1c73e697;
assign   tb_o_tag_ready[637]                  =   1'b0;
assign   tb_o_tag[637]                        =   tb_o_tag[636];

// CLK no. 638/1240
// *************************************************
assign   tb_i_valid[638]                      =   1'b0;
assign   tb_i_reset[638]                      =   1'b0;
assign   tb_i_sop[638]                        =   1'b0;
assign   tb_i_key_update[638]                 =   1'b0;
assign   tb_i_key[638]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[638]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[638]               =   1'b0;
assign   tb_i_rf_static_encrypt[638]          =   1'b1;
assign   tb_i_clear_fault_flags[638]          =   1'b0;
assign   tb_i_rf_static_aad_length[638]       =   64'h0000000000000100;
assign   tb_i_aad[638]                        =   tb_i_aad[637];
assign   tb_i_rf_static_plaintext_length[638] =   64'h0000000000000280;
assign   tb_i_plaintext[638]                  =   tb_i_plaintext[637];
assign   tb_o_valid[638]                      =   1'b1;
assign   tb_o_sop[638]                        =   1'b0;
assign   tb_o_ciphertext[638]                 =   256'hb7cf748c22cd87d749ed3a64e7d0f9b02e32910a36b242182c00e4c826ab60bf;
assign   tb_o_tag_ready[638]                  =   1'b0;
assign   tb_o_tag[638]                        =   tb_o_tag[637];

// CLK no. 639/1240
// *************************************************
assign   tb_i_valid[639]                      =   1'b0;
assign   tb_i_reset[639]                      =   1'b0;
assign   tb_i_sop[639]                        =   1'b0;
assign   tb_i_key_update[639]                 =   1'b0;
assign   tb_i_key[639]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[639]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[639]               =   1'b0;
assign   tb_i_rf_static_encrypt[639]          =   1'b1;
assign   tb_i_clear_fault_flags[639]          =   1'b0;
assign   tb_i_rf_static_aad_length[639]       =   64'h0000000000000100;
assign   tb_i_aad[639]                        =   tb_i_aad[638];
assign   tb_i_rf_static_plaintext_length[639] =   64'h0000000000000280;
assign   tb_i_plaintext[639]                  =   tb_i_plaintext[638];
assign   tb_o_valid[639]                      =   1'b1;
assign   tb_o_sop[639]                        =   1'b0;
assign   tb_o_ciphertext[639]                 =   256'h883e9351111aa2c93ab17905c35615f6;
assign   tb_o_tag_ready[639]                  =   1'b0;
assign   tb_o_tag[639]                        =   tb_o_tag[638];

// CLK no. 640/1240
// *************************************************
assign   tb_i_valid[640]                      =   1'b0;
assign   tb_i_reset[640]                      =   1'b0;
assign   tb_i_sop[640]                        =   1'b0;
assign   tb_i_key_update[640]                 =   1'b0;
assign   tb_i_key[640]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[640]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[640]               =   1'b0;
assign   tb_i_rf_static_encrypt[640]          =   1'b1;
assign   tb_i_clear_fault_flags[640]          =   1'b0;
assign   tb_i_rf_static_aad_length[640]       =   64'h0000000000000100;
assign   tb_i_aad[640]                        =   tb_i_aad[639];
assign   tb_i_rf_static_plaintext_length[640] =   64'h0000000000000280;
assign   tb_i_plaintext[640]                  =   tb_i_plaintext[639];
assign   tb_o_valid[640]                      =   1'b0;
assign   tb_o_sop[640]                        =   1'b0;
assign   tb_o_ciphertext[640]                 =   tb_o_ciphertext[639];
assign   tb_o_tag_ready[640]                  =   1'b0;
assign   tb_o_tag[640]                        =   tb_o_tag[639];

// CLK no. 641/1240
// *************************************************
assign   tb_i_valid[641]                      =   1'b0;
assign   tb_i_reset[641]                      =   1'b0;
assign   tb_i_sop[641]                        =   1'b0;
assign   tb_i_key_update[641]                 =   1'b0;
assign   tb_i_key[641]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[641]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[641]               =   1'b0;
assign   tb_i_rf_static_encrypt[641]          =   1'b1;
assign   tb_i_clear_fault_flags[641]          =   1'b0;
assign   tb_i_rf_static_aad_length[641]       =   64'h0000000000000100;
assign   tb_i_aad[641]                        =   tb_i_aad[640];
assign   tb_i_rf_static_plaintext_length[641] =   64'h0000000000000280;
assign   tb_i_plaintext[641]                  =   tb_i_plaintext[640];
assign   tb_o_valid[641]                      =   1'b0;
assign   tb_o_sop[641]                        =   1'b0;
assign   tb_o_ciphertext[641]                 =   tb_o_ciphertext[640];
assign   tb_o_tag_ready[641]                  =   1'b0;
assign   tb_o_tag[641]                        =   tb_o_tag[640];

// CLK no. 642/1240
// *************************************************
assign   tb_i_valid[642]                      =   1'b0;
assign   tb_i_reset[642]                      =   1'b0;
assign   tb_i_sop[642]                        =   1'b0;
assign   tb_i_key_update[642]                 =   1'b0;
assign   tb_i_key[642]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[642]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[642]               =   1'b0;
assign   tb_i_rf_static_encrypt[642]          =   1'b1;
assign   tb_i_clear_fault_flags[642]          =   1'b0;
assign   tb_i_rf_static_aad_length[642]       =   64'h0000000000000100;
assign   tb_i_aad[642]                        =   tb_i_aad[641];
assign   tb_i_rf_static_plaintext_length[642] =   64'h0000000000000280;
assign   tb_i_plaintext[642]                  =   tb_i_plaintext[641];
assign   tb_o_valid[642]                      =   1'b0;
assign   tb_o_sop[642]                        =   1'b0;
assign   tb_o_ciphertext[642]                 =   tb_o_ciphertext[641];
assign   tb_o_tag_ready[642]                  =   1'b0;
assign   tb_o_tag[642]                        =   tb_o_tag[641];

// CLK no. 643/1240
// *************************************************
assign   tb_i_valid[643]                      =   1'b0;
assign   tb_i_reset[643]                      =   1'b0;
assign   tb_i_sop[643]                        =   1'b0;
assign   tb_i_key_update[643]                 =   1'b0;
assign   tb_i_key[643]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[643]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[643]               =   1'b0;
assign   tb_i_rf_static_encrypt[643]          =   1'b1;
assign   tb_i_clear_fault_flags[643]          =   1'b0;
assign   tb_i_rf_static_aad_length[643]       =   64'h0000000000000100;
assign   tb_i_aad[643]                        =   tb_i_aad[642];
assign   tb_i_rf_static_plaintext_length[643] =   64'h0000000000000280;
assign   tb_i_plaintext[643]                  =   tb_i_plaintext[642];
assign   tb_o_valid[643]                      =   1'b0;
assign   tb_o_sop[643]                        =   1'b0;
assign   tb_o_ciphertext[643]                 =   tb_o_ciphertext[642];
assign   tb_o_tag_ready[643]                  =   1'b0;
assign   tb_o_tag[643]                        =   tb_o_tag[642];

// CLK no. 644/1240
// *************************************************
assign   tb_i_valid[644]                      =   1'b0;
assign   tb_i_reset[644]                      =   1'b0;
assign   tb_i_sop[644]                        =   1'b0;
assign   tb_i_key_update[644]                 =   1'b0;
assign   tb_i_key[644]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[644]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[644]               =   1'b0;
assign   tb_i_rf_static_encrypt[644]          =   1'b1;
assign   tb_i_clear_fault_flags[644]          =   1'b0;
assign   tb_i_rf_static_aad_length[644]       =   64'h0000000000000100;
assign   tb_i_aad[644]                        =   tb_i_aad[643];
assign   tb_i_rf_static_plaintext_length[644] =   64'h0000000000000280;
assign   tb_i_plaintext[644]                  =   tb_i_plaintext[643];
assign   tb_o_valid[644]                      =   1'b0;
assign   tb_o_sop[644]                        =   1'b0;
assign   tb_o_ciphertext[644]                 =   tb_o_ciphertext[643];
assign   tb_o_tag_ready[644]                  =   1'b0;
assign   tb_o_tag[644]                        =   tb_o_tag[643];

// CLK no. 645/1240
// *************************************************
assign   tb_i_valid[645]                      =   1'b0;
assign   tb_i_reset[645]                      =   1'b0;
assign   tb_i_sop[645]                        =   1'b0;
assign   tb_i_key_update[645]                 =   1'b0;
assign   tb_i_key[645]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[645]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[645]               =   1'b0;
assign   tb_i_rf_static_encrypt[645]          =   1'b1;
assign   tb_i_clear_fault_flags[645]          =   1'b0;
assign   tb_i_rf_static_aad_length[645]       =   64'h0000000000000100;
assign   tb_i_aad[645]                        =   tb_i_aad[644];
assign   tb_i_rf_static_plaintext_length[645] =   64'h0000000000000280;
assign   tb_i_plaintext[645]                  =   tb_i_plaintext[644];
assign   tb_o_valid[645]                      =   1'b0;
assign   tb_o_sop[645]                        =   1'b0;
assign   tb_o_ciphertext[645]                 =   tb_o_ciphertext[644];
assign   tb_o_tag_ready[645]                  =   1'b0;
assign   tb_o_tag[645]                        =   tb_o_tag[644];

// CLK no. 646/1240
// *************************************************
assign   tb_i_valid[646]                      =   1'b0;
assign   tb_i_reset[646]                      =   1'b0;
assign   tb_i_sop[646]                        =   1'b0;
assign   tb_i_key_update[646]                 =   1'b0;
assign   tb_i_key[646]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[646]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[646]               =   1'b0;
assign   tb_i_rf_static_encrypt[646]          =   1'b1;
assign   tb_i_clear_fault_flags[646]          =   1'b0;
assign   tb_i_rf_static_aad_length[646]       =   64'h0000000000000100;
assign   tb_i_aad[646]                        =   tb_i_aad[645];
assign   tb_i_rf_static_plaintext_length[646] =   64'h0000000000000280;
assign   tb_i_plaintext[646]                  =   tb_i_plaintext[645];
assign   tb_o_valid[646]                      =   1'b0;
assign   tb_o_sop[646]                        =   1'b0;
assign   tb_o_ciphertext[646]                 =   tb_o_ciphertext[645];
assign   tb_o_tag_ready[646]                  =   1'b0;
assign   tb_o_tag[646]                        =   tb_o_tag[645];

// CLK no. 647/1240
// *************************************************
assign   tb_i_valid[647]                      =   1'b0;
assign   tb_i_reset[647]                      =   1'b0;
assign   tb_i_sop[647]                        =   1'b0;
assign   tb_i_key_update[647]                 =   1'b0;
assign   tb_i_key[647]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[647]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[647]               =   1'b0;
assign   tb_i_rf_static_encrypt[647]          =   1'b1;
assign   tb_i_clear_fault_flags[647]          =   1'b0;
assign   tb_i_rf_static_aad_length[647]       =   64'h0000000000000100;
assign   tb_i_aad[647]                        =   tb_i_aad[646];
assign   tb_i_rf_static_plaintext_length[647] =   64'h0000000000000280;
assign   tb_i_plaintext[647]                  =   tb_i_plaintext[646];
assign   tb_o_valid[647]                      =   1'b0;
assign   tb_o_sop[647]                        =   1'b0;
assign   tb_o_ciphertext[647]                 =   tb_o_ciphertext[646];
assign   tb_o_tag_ready[647]                  =   1'b1;
assign   tb_o_tag[647]                        =   128'h70943eca1e63481cf3c561084722bdf7;

// CLK no. 648/1240
// *************************************************
assign   tb_i_valid[648]                      =   1'b0;
assign   tb_i_reset[648]                      =   1'b0;
assign   tb_i_sop[648]                        =   1'b0;
assign   tb_i_key_update[648]                 =   1'b0;
assign   tb_i_key[648]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[648]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[648]               =   1'b0;
assign   tb_i_rf_static_encrypt[648]          =   1'b1;
assign   tb_i_clear_fault_flags[648]          =   1'b0;
assign   tb_i_rf_static_aad_length[648]       =   64'h0000000000000100;
assign   tb_i_aad[648]                        =   tb_i_aad[647];
assign   tb_i_rf_static_plaintext_length[648] =   64'h0000000000000280;
assign   tb_i_plaintext[648]                  =   tb_i_plaintext[647];
assign   tb_o_valid[648]                      =   1'b0;
assign   tb_o_sop[648]                        =   1'b0;
assign   tb_o_ciphertext[648]                 =   tb_o_ciphertext[647];
assign   tb_o_tag_ready[648]                  =   1'b0;
assign   tb_o_tag[648]                        =   tb_o_tag[647];

// CLK no. 649/1240
// *************************************************
assign   tb_i_valid[649]                      =   1'b0;
assign   tb_i_reset[649]                      =   1'b0;
assign   tb_i_sop[649]                        =   1'b0;
assign   tb_i_key_update[649]                 =   1'b0;
assign   tb_i_key[649]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[649]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[649]               =   1'b0;
assign   tb_i_rf_static_encrypt[649]          =   1'b1;
assign   tb_i_clear_fault_flags[649]          =   1'b0;
assign   tb_i_rf_static_aad_length[649]       =   64'h0000000000000100;
assign   tb_i_aad[649]                        =   tb_i_aad[648];
assign   tb_i_rf_static_plaintext_length[649] =   64'h0000000000000280;
assign   tb_i_plaintext[649]                  =   tb_i_plaintext[648];
assign   tb_o_valid[649]                      =   1'b0;
assign   tb_o_sop[649]                        =   1'b0;
assign   tb_o_ciphertext[649]                 =   tb_o_ciphertext[648];
assign   tb_o_tag_ready[649]                  =   1'b0;
assign   tb_o_tag[649]                        =   tb_o_tag[648];

// CLK no. 650/1240
// *************************************************
assign   tb_i_valid[650]                      =   1'b0;
assign   tb_i_reset[650]                      =   1'b0;
assign   tb_i_sop[650]                        =   1'b1;
assign   tb_i_key_update[650]                 =   1'b0;
assign   tb_i_key[650]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[650]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[650]               =   1'b0;
assign   tb_i_rf_static_encrypt[650]          =   1'b1;
assign   tb_i_clear_fault_flags[650]          =   1'b0;
assign   tb_i_rf_static_aad_length[650]       =   64'h0000000000000100;
assign   tb_i_aad[650]                        =   tb_i_aad[649];
assign   tb_i_rf_static_plaintext_length[650] =   64'h0000000000000280;
assign   tb_i_plaintext[650]                  =   tb_i_plaintext[649];
assign   tb_o_valid[650]                      =   1'b0;
assign   tb_o_sop[650]                        =   1'b0;
assign   tb_o_ciphertext[650]                 =   tb_o_ciphertext[649];
assign   tb_o_tag_ready[650]                  =   1'b0;
assign   tb_o_tag[650]                        =   tb_o_tag[649];

// CLK no. 651/1240
// *************************************************
assign   tb_i_valid[651]                      =   1'b1;
assign   tb_i_reset[651]                      =   1'b0;
assign   tb_i_sop[651]                        =   1'b0;
assign   tb_i_key_update[651]                 =   1'b0;
assign   tb_i_key[651]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[651]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[651]               =   1'b0;
assign   tb_i_rf_static_encrypt[651]          =   1'b1;
assign   tb_i_clear_fault_flags[651]          =   1'b0;
assign   tb_i_rf_static_aad_length[651]       =   64'h0000000000000100;
assign   tb_i_aad[651]                        =   256'h21beb7686494ef29dba2fd29183b28441723ca31397d67dcd3ee879e6b2fb488;
assign   tb_i_rf_static_plaintext_length[651] =   64'h0000000000000280;
assign   tb_i_plaintext[651]                  =   tb_i_plaintext[650];
assign   tb_o_valid[651]                      =   1'b0;
assign   tb_o_sop[651]                        =   1'b0;
assign   tb_o_ciphertext[651]                 =   tb_o_ciphertext[650];
assign   tb_o_tag_ready[651]                  =   1'b0;
assign   tb_o_tag[651]                        =   tb_o_tag[650];

// CLK no. 652/1240
// *************************************************
assign   tb_i_valid[652]                      =   1'b1;
assign   tb_i_reset[652]                      =   1'b0;
assign   tb_i_sop[652]                        =   1'b0;
assign   tb_i_key_update[652]                 =   1'b0;
assign   tb_i_key[652]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[652]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[652]               =   1'b0;
assign   tb_i_rf_static_encrypt[652]          =   1'b1;
assign   tb_i_clear_fault_flags[652]          =   1'b0;
assign   tb_i_rf_static_aad_length[652]       =   64'h0000000000000100;
assign   tb_i_aad[652]                        =   tb_i_aad[651];
assign   tb_i_rf_static_plaintext_length[652] =   64'h0000000000000280;
assign   tb_i_plaintext[652]                  =   256'hbdf1adfb6ce61887fce2397e217ce90ceaeb197a9eb36a2d87648350439f2fda;
assign   tb_o_valid[652]                      =   1'b0;
assign   tb_o_sop[652]                        =   1'b0;
assign   tb_o_ciphertext[652]                 =   tb_o_ciphertext[651];
assign   tb_o_tag_ready[652]                  =   1'b0;
assign   tb_o_tag[652]                        =   tb_o_tag[651];

// CLK no. 653/1240
// *************************************************
assign   tb_i_valid[653]                      =   1'b1;
assign   tb_i_reset[653]                      =   1'b0;
assign   tb_i_sop[653]                        =   1'b0;
assign   tb_i_key_update[653]                 =   1'b0;
assign   tb_i_key[653]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[653]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[653]               =   1'b0;
assign   tb_i_rf_static_encrypt[653]          =   1'b1;
assign   tb_i_clear_fault_flags[653]          =   1'b0;
assign   tb_i_rf_static_aad_length[653]       =   64'h0000000000000100;
assign   tb_i_aad[653]                        =   tb_i_aad[652];
assign   tb_i_rf_static_plaintext_length[653] =   64'h0000000000000280;
assign   tb_i_plaintext[653]                  =   256'hfdbb556c6a2278ccb69cafbd25e1cfbe4cd7f14f50451bc54ff34cf7c2fedd03;
assign   tb_o_valid[653]                      =   1'b0;
assign   tb_o_sop[653]                        =   1'b0;
assign   tb_o_ciphertext[653]                 =   tb_o_ciphertext[652];
assign   tb_o_tag_ready[653]                  =   1'b0;
assign   tb_o_tag[653]                        =   tb_o_tag[652];

// CLK no. 654/1240
// *************************************************
assign   tb_i_valid[654]                      =   1'b1;
assign   tb_i_reset[654]                      =   1'b0;
assign   tb_i_sop[654]                        =   1'b0;
assign   tb_i_key_update[654]                 =   1'b0;
assign   tb_i_key[654]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[654]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[654]               =   1'b0;
assign   tb_i_rf_static_encrypt[654]          =   1'b1;
assign   tb_i_clear_fault_flags[654]          =   1'b0;
assign   tb_i_rf_static_aad_length[654]       =   64'h0000000000000100;
assign   tb_i_aad[654]                        =   tb_i_aad[653];
assign   tb_i_rf_static_plaintext_length[654] =   64'h0000000000000280;
assign   tb_i_plaintext[654]                  =   256'hdf617264153455d39da68bc1cd574117;
assign   tb_o_valid[654]                      =   1'b0;
assign   tb_o_sop[654]                        =   1'b0;
assign   tb_o_ciphertext[654]                 =   tb_o_ciphertext[653];
assign   tb_o_tag_ready[654]                  =   1'b0;
assign   tb_o_tag[654]                        =   tb_o_tag[653];

// CLK no. 655/1240
// *************************************************
assign   tb_i_valid[655]                      =   1'b0;
assign   tb_i_reset[655]                      =   1'b0;
assign   tb_i_sop[655]                        =   1'b0;
assign   tb_i_key_update[655]                 =   1'b0;
assign   tb_i_key[655]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[655]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[655]               =   1'b0;
assign   tb_i_rf_static_encrypt[655]          =   1'b1;
assign   tb_i_clear_fault_flags[655]          =   1'b0;
assign   tb_i_rf_static_aad_length[655]       =   64'h0000000000000100;
assign   tb_i_aad[655]                        =   tb_i_aad[654];
assign   tb_i_rf_static_plaintext_length[655] =   64'h0000000000000280;
assign   tb_i_plaintext[655]                  =   tb_i_plaintext[654];
assign   tb_o_valid[655]                      =   1'b0;
assign   tb_o_sop[655]                        =   1'b0;
assign   tb_o_ciphertext[655]                 =   tb_o_ciphertext[654];
assign   tb_o_tag_ready[655]                  =   1'b0;
assign   tb_o_tag[655]                        =   tb_o_tag[654];

// CLK no. 656/1240
// *************************************************
assign   tb_i_valid[656]                      =   1'b0;
assign   tb_i_reset[656]                      =   1'b0;
assign   tb_i_sop[656]                        =   1'b0;
assign   tb_i_key_update[656]                 =   1'b0;
assign   tb_i_key[656]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[656]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[656]               =   1'b0;
assign   tb_i_rf_static_encrypt[656]          =   1'b1;
assign   tb_i_clear_fault_flags[656]          =   1'b0;
assign   tb_i_rf_static_aad_length[656]       =   64'h0000000000000100;
assign   tb_i_aad[656]                        =   tb_i_aad[655];
assign   tb_i_rf_static_plaintext_length[656] =   64'h0000000000000280;
assign   tb_i_plaintext[656]                  =   tb_i_plaintext[655];
assign   tb_o_valid[656]                      =   1'b0;
assign   tb_o_sop[656]                        =   1'b0;
assign   tb_o_ciphertext[656]                 =   tb_o_ciphertext[655];
assign   tb_o_tag_ready[656]                  =   1'b0;
assign   tb_o_tag[656]                        =   tb_o_tag[655];

// CLK no. 657/1240
// *************************************************
assign   tb_i_valid[657]                      =   1'b0;
assign   tb_i_reset[657]                      =   1'b0;
assign   tb_i_sop[657]                        =   1'b0;
assign   tb_i_key_update[657]                 =   1'b0;
assign   tb_i_key[657]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[657]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[657]               =   1'b0;
assign   tb_i_rf_static_encrypt[657]          =   1'b1;
assign   tb_i_clear_fault_flags[657]          =   1'b0;
assign   tb_i_rf_static_aad_length[657]       =   64'h0000000000000100;
assign   tb_i_aad[657]                        =   tb_i_aad[656];
assign   tb_i_rf_static_plaintext_length[657] =   64'h0000000000000280;
assign   tb_i_plaintext[657]                  =   tb_i_plaintext[656];
assign   tb_o_valid[657]                      =   1'b0;
assign   tb_o_sop[657]                        =   1'b0;
assign   tb_o_ciphertext[657]                 =   tb_o_ciphertext[656];
assign   tb_o_tag_ready[657]                  =   1'b0;
assign   tb_o_tag[657]                        =   tb_o_tag[656];

// CLK no. 658/1240
// *************************************************
assign   tb_i_valid[658]                      =   1'b0;
assign   tb_i_reset[658]                      =   1'b0;
assign   tb_i_sop[658]                        =   1'b0;
assign   tb_i_key_update[658]                 =   1'b0;
assign   tb_i_key[658]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[658]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[658]               =   1'b0;
assign   tb_i_rf_static_encrypt[658]          =   1'b1;
assign   tb_i_clear_fault_flags[658]          =   1'b0;
assign   tb_i_rf_static_aad_length[658]       =   64'h0000000000000100;
assign   tb_i_aad[658]                        =   tb_i_aad[657];
assign   tb_i_rf_static_plaintext_length[658] =   64'h0000000000000280;
assign   tb_i_plaintext[658]                  =   tb_i_plaintext[657];
assign   tb_o_valid[658]                      =   1'b0;
assign   tb_o_sop[658]                        =   1'b0;
assign   tb_o_ciphertext[658]                 =   tb_o_ciphertext[657];
assign   tb_o_tag_ready[658]                  =   1'b0;
assign   tb_o_tag[658]                        =   tb_o_tag[657];

// CLK no. 659/1240
// *************************************************
assign   tb_i_valid[659]                      =   1'b0;
assign   tb_i_reset[659]                      =   1'b0;
assign   tb_i_sop[659]                        =   1'b0;
assign   tb_i_key_update[659]                 =   1'b0;
assign   tb_i_key[659]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[659]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[659]               =   1'b0;
assign   tb_i_rf_static_encrypt[659]          =   1'b1;
assign   tb_i_clear_fault_flags[659]          =   1'b0;
assign   tb_i_rf_static_aad_length[659]       =   64'h0000000000000100;
assign   tb_i_aad[659]                        =   tb_i_aad[658];
assign   tb_i_rf_static_plaintext_length[659] =   64'h0000000000000280;
assign   tb_i_plaintext[659]                  =   tb_i_plaintext[658];
assign   tb_o_valid[659]                      =   1'b0;
assign   tb_o_sop[659]                        =   1'b0;
assign   tb_o_ciphertext[659]                 =   tb_o_ciphertext[658];
assign   tb_o_tag_ready[659]                  =   1'b0;
assign   tb_o_tag[659]                        =   tb_o_tag[658];

// CLK no. 660/1240
// *************************************************
assign   tb_i_valid[660]                      =   1'b0;
assign   tb_i_reset[660]                      =   1'b0;
assign   tb_i_sop[660]                        =   1'b0;
assign   tb_i_key_update[660]                 =   1'b0;
assign   tb_i_key[660]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[660]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[660]               =   1'b0;
assign   tb_i_rf_static_encrypt[660]          =   1'b1;
assign   tb_i_clear_fault_flags[660]          =   1'b0;
assign   tb_i_rf_static_aad_length[660]       =   64'h0000000000000100;
assign   tb_i_aad[660]                        =   tb_i_aad[659];
assign   tb_i_rf_static_plaintext_length[660] =   64'h0000000000000280;
assign   tb_i_plaintext[660]                  =   tb_i_plaintext[659];
assign   tb_o_valid[660]                      =   1'b0;
assign   tb_o_sop[660]                        =   1'b0;
assign   tb_o_ciphertext[660]                 =   tb_o_ciphertext[659];
assign   tb_o_tag_ready[660]                  =   1'b0;
assign   tb_o_tag[660]                        =   tb_o_tag[659];

// CLK no. 661/1240
// *************************************************
assign   tb_i_valid[661]                      =   1'b0;
assign   tb_i_reset[661]                      =   1'b0;
assign   tb_i_sop[661]                        =   1'b0;
assign   tb_i_key_update[661]                 =   1'b0;
assign   tb_i_key[661]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[661]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[661]               =   1'b0;
assign   tb_i_rf_static_encrypt[661]          =   1'b1;
assign   tb_i_clear_fault_flags[661]          =   1'b0;
assign   tb_i_rf_static_aad_length[661]       =   64'h0000000000000100;
assign   tb_i_aad[661]                        =   tb_i_aad[660];
assign   tb_i_rf_static_plaintext_length[661] =   64'h0000000000000280;
assign   tb_i_plaintext[661]                  =   tb_i_plaintext[660];
assign   tb_o_valid[661]                      =   1'b0;
assign   tb_o_sop[661]                        =   1'b0;
assign   tb_o_ciphertext[661]                 =   tb_o_ciphertext[660];
assign   tb_o_tag_ready[661]                  =   1'b0;
assign   tb_o_tag[661]                        =   tb_o_tag[660];

// CLK no. 662/1240
// *************************************************
assign   tb_i_valid[662]                      =   1'b0;
assign   tb_i_reset[662]                      =   1'b0;
assign   tb_i_sop[662]                        =   1'b0;
assign   tb_i_key_update[662]                 =   1'b0;
assign   tb_i_key[662]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[662]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[662]               =   1'b0;
assign   tb_i_rf_static_encrypt[662]          =   1'b1;
assign   tb_i_clear_fault_flags[662]          =   1'b0;
assign   tb_i_rf_static_aad_length[662]       =   64'h0000000000000100;
assign   tb_i_aad[662]                        =   tb_i_aad[661];
assign   tb_i_rf_static_plaintext_length[662] =   64'h0000000000000280;
assign   tb_i_plaintext[662]                  =   tb_i_plaintext[661];
assign   tb_o_valid[662]                      =   1'b0;
assign   tb_o_sop[662]                        =   1'b0;
assign   tb_o_ciphertext[662]                 =   tb_o_ciphertext[661];
assign   tb_o_tag_ready[662]                  =   1'b0;
assign   tb_o_tag[662]                        =   tb_o_tag[661];

// CLK no. 663/1240
// *************************************************
assign   tb_i_valid[663]                      =   1'b0;
assign   tb_i_reset[663]                      =   1'b0;
assign   tb_i_sop[663]                        =   1'b0;
assign   tb_i_key_update[663]                 =   1'b0;
assign   tb_i_key[663]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[663]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[663]               =   1'b0;
assign   tb_i_rf_static_encrypt[663]          =   1'b1;
assign   tb_i_clear_fault_flags[663]          =   1'b0;
assign   tb_i_rf_static_aad_length[663]       =   64'h0000000000000100;
assign   tb_i_aad[663]                        =   tb_i_aad[662];
assign   tb_i_rf_static_plaintext_length[663] =   64'h0000000000000280;
assign   tb_i_plaintext[663]                  =   tb_i_plaintext[662];
assign   tb_o_valid[663]                      =   1'b0;
assign   tb_o_sop[663]                        =   1'b0;
assign   tb_o_ciphertext[663]                 =   tb_o_ciphertext[662];
assign   tb_o_tag_ready[663]                  =   1'b0;
assign   tb_o_tag[663]                        =   tb_o_tag[662];

// CLK no. 664/1240
// *************************************************
assign   tb_i_valid[664]                      =   1'b0;
assign   tb_i_reset[664]                      =   1'b0;
assign   tb_i_sop[664]                        =   1'b0;
assign   tb_i_key_update[664]                 =   1'b0;
assign   tb_i_key[664]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[664]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[664]               =   1'b0;
assign   tb_i_rf_static_encrypt[664]          =   1'b1;
assign   tb_i_clear_fault_flags[664]          =   1'b0;
assign   tb_i_rf_static_aad_length[664]       =   64'h0000000000000100;
assign   tb_i_aad[664]                        =   tb_i_aad[663];
assign   tb_i_rf_static_plaintext_length[664] =   64'h0000000000000280;
assign   tb_i_plaintext[664]                  =   tb_i_plaintext[663];
assign   tb_o_valid[664]                      =   1'b0;
assign   tb_o_sop[664]                        =   1'b0;
assign   tb_o_ciphertext[664]                 =   tb_o_ciphertext[663];
assign   tb_o_tag_ready[664]                  =   1'b0;
assign   tb_o_tag[664]                        =   tb_o_tag[663];

// CLK no. 665/1240
// *************************************************
assign   tb_i_valid[665]                      =   1'b0;
assign   tb_i_reset[665]                      =   1'b0;
assign   tb_i_sop[665]                        =   1'b0;
assign   tb_i_key_update[665]                 =   1'b0;
assign   tb_i_key[665]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[665]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[665]               =   1'b0;
assign   tb_i_rf_static_encrypt[665]          =   1'b1;
assign   tb_i_clear_fault_flags[665]          =   1'b0;
assign   tb_i_rf_static_aad_length[665]       =   64'h0000000000000100;
assign   tb_i_aad[665]                        =   tb_i_aad[664];
assign   tb_i_rf_static_plaintext_length[665] =   64'h0000000000000280;
assign   tb_i_plaintext[665]                  =   tb_i_plaintext[664];
assign   tb_o_valid[665]                      =   1'b0;
assign   tb_o_sop[665]                        =   1'b0;
assign   tb_o_ciphertext[665]                 =   tb_o_ciphertext[664];
assign   tb_o_tag_ready[665]                  =   1'b0;
assign   tb_o_tag[665]                        =   tb_o_tag[664];

// CLK no. 666/1240
// *************************************************
assign   tb_i_valid[666]                      =   1'b0;
assign   tb_i_reset[666]                      =   1'b0;
assign   tb_i_sop[666]                        =   1'b0;
assign   tb_i_key_update[666]                 =   1'b0;
assign   tb_i_key[666]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[666]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[666]               =   1'b0;
assign   tb_i_rf_static_encrypt[666]          =   1'b1;
assign   tb_i_clear_fault_flags[666]          =   1'b0;
assign   tb_i_rf_static_aad_length[666]       =   64'h0000000000000100;
assign   tb_i_aad[666]                        =   tb_i_aad[665];
assign   tb_i_rf_static_plaintext_length[666] =   64'h0000000000000280;
assign   tb_i_plaintext[666]                  =   tb_i_plaintext[665];
assign   tb_o_valid[666]                      =   1'b0;
assign   tb_o_sop[666]                        =   1'b0;
assign   tb_o_ciphertext[666]                 =   tb_o_ciphertext[665];
assign   tb_o_tag_ready[666]                  =   1'b0;
assign   tb_o_tag[666]                        =   tb_o_tag[665];

// CLK no. 667/1240
// *************************************************
assign   tb_i_valid[667]                      =   1'b0;
assign   tb_i_reset[667]                      =   1'b0;
assign   tb_i_sop[667]                        =   1'b0;
assign   tb_i_key_update[667]                 =   1'b0;
assign   tb_i_key[667]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[667]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[667]               =   1'b0;
assign   tb_i_rf_static_encrypt[667]          =   1'b1;
assign   tb_i_clear_fault_flags[667]          =   1'b0;
assign   tb_i_rf_static_aad_length[667]       =   64'h0000000000000100;
assign   tb_i_aad[667]                        =   tb_i_aad[666];
assign   tb_i_rf_static_plaintext_length[667] =   64'h0000000000000280;
assign   tb_i_plaintext[667]                  =   tb_i_plaintext[666];
assign   tb_o_valid[667]                      =   1'b0;
assign   tb_o_sop[667]                        =   1'b0;
assign   tb_o_ciphertext[667]                 =   tb_o_ciphertext[666];
assign   tb_o_tag_ready[667]                  =   1'b0;
assign   tb_o_tag[667]                        =   tb_o_tag[666];

// CLK no. 668/1240
// *************************************************
assign   tb_i_valid[668]                      =   1'b0;
assign   tb_i_reset[668]                      =   1'b0;
assign   tb_i_sop[668]                        =   1'b0;
assign   tb_i_key_update[668]                 =   1'b0;
assign   tb_i_key[668]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[668]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[668]               =   1'b0;
assign   tb_i_rf_static_encrypt[668]          =   1'b1;
assign   tb_i_clear_fault_flags[668]          =   1'b0;
assign   tb_i_rf_static_aad_length[668]       =   64'h0000000000000100;
assign   tb_i_aad[668]                        =   tb_i_aad[667];
assign   tb_i_rf_static_plaintext_length[668] =   64'h0000000000000280;
assign   tb_i_plaintext[668]                  =   tb_i_plaintext[667];
assign   tb_o_valid[668]                      =   1'b0;
assign   tb_o_sop[668]                        =   1'b0;
assign   tb_o_ciphertext[668]                 =   tb_o_ciphertext[667];
assign   tb_o_tag_ready[668]                  =   1'b0;
assign   tb_o_tag[668]                        =   tb_o_tag[667];

// CLK no. 669/1240
// *************************************************
assign   tb_i_valid[669]                      =   1'b0;
assign   tb_i_reset[669]                      =   1'b0;
assign   tb_i_sop[669]                        =   1'b0;
assign   tb_i_key_update[669]                 =   1'b0;
assign   tb_i_key[669]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[669]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[669]               =   1'b0;
assign   tb_i_rf_static_encrypt[669]          =   1'b1;
assign   tb_i_clear_fault_flags[669]          =   1'b0;
assign   tb_i_rf_static_aad_length[669]       =   64'h0000000000000100;
assign   tb_i_aad[669]                        =   tb_i_aad[668];
assign   tb_i_rf_static_plaintext_length[669] =   64'h0000000000000280;
assign   tb_i_plaintext[669]                  =   tb_i_plaintext[668];
assign   tb_o_valid[669]                      =   1'b0;
assign   tb_o_sop[669]                        =   1'b0;
assign   tb_o_ciphertext[669]                 =   tb_o_ciphertext[668];
assign   tb_o_tag_ready[669]                  =   1'b0;
assign   tb_o_tag[669]                        =   tb_o_tag[668];

// CLK no. 670/1240
// *************************************************
assign   tb_i_valid[670]                      =   1'b0;
assign   tb_i_reset[670]                      =   1'b0;
assign   tb_i_sop[670]                        =   1'b0;
assign   tb_i_key_update[670]                 =   1'b0;
assign   tb_i_key[670]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[670]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[670]               =   1'b0;
assign   tb_i_rf_static_encrypt[670]          =   1'b1;
assign   tb_i_clear_fault_flags[670]          =   1'b0;
assign   tb_i_rf_static_aad_length[670]       =   64'h0000000000000100;
assign   tb_i_aad[670]                        =   tb_i_aad[669];
assign   tb_i_rf_static_plaintext_length[670] =   64'h0000000000000280;
assign   tb_i_plaintext[670]                  =   tb_i_plaintext[669];
assign   tb_o_valid[670]                      =   1'b0;
assign   tb_o_sop[670]                        =   1'b0;
assign   tb_o_ciphertext[670]                 =   tb_o_ciphertext[669];
assign   tb_o_tag_ready[670]                  =   1'b0;
assign   tb_o_tag[670]                        =   tb_o_tag[669];

// CLK no. 671/1240
// *************************************************
assign   tb_i_valid[671]                      =   1'b0;
assign   tb_i_reset[671]                      =   1'b0;
assign   tb_i_sop[671]                        =   1'b0;
assign   tb_i_key_update[671]                 =   1'b0;
assign   tb_i_key[671]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[671]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[671]               =   1'b0;
assign   tb_i_rf_static_encrypt[671]          =   1'b1;
assign   tb_i_clear_fault_flags[671]          =   1'b0;
assign   tb_i_rf_static_aad_length[671]       =   64'h0000000000000100;
assign   tb_i_aad[671]                        =   tb_i_aad[670];
assign   tb_i_rf_static_plaintext_length[671] =   64'h0000000000000280;
assign   tb_i_plaintext[671]                  =   tb_i_plaintext[670];
assign   tb_o_valid[671]                      =   1'b0;
assign   tb_o_sop[671]                        =   1'b0;
assign   tb_o_ciphertext[671]                 =   tb_o_ciphertext[670];
assign   tb_o_tag_ready[671]                  =   1'b0;
assign   tb_o_tag[671]                        =   tb_o_tag[670];

// CLK no. 672/1240
// *************************************************
assign   tb_i_valid[672]                      =   1'b0;
assign   tb_i_reset[672]                      =   1'b0;
assign   tb_i_sop[672]                        =   1'b0;
assign   tb_i_key_update[672]                 =   1'b0;
assign   tb_i_key[672]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[672]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[672]               =   1'b0;
assign   tb_i_rf_static_encrypt[672]          =   1'b1;
assign   tb_i_clear_fault_flags[672]          =   1'b0;
assign   tb_i_rf_static_aad_length[672]       =   64'h0000000000000100;
assign   tb_i_aad[672]                        =   tb_i_aad[671];
assign   tb_i_rf_static_plaintext_length[672] =   64'h0000000000000280;
assign   tb_i_plaintext[672]                  =   tb_i_plaintext[671];
assign   tb_o_valid[672]                      =   1'b0;
assign   tb_o_sop[672]                        =   1'b0;
assign   tb_o_ciphertext[672]                 =   tb_o_ciphertext[671];
assign   tb_o_tag_ready[672]                  =   1'b0;
assign   tb_o_tag[672]                        =   tb_o_tag[671];

// CLK no. 673/1240
// *************************************************
assign   tb_i_valid[673]                      =   1'b0;
assign   tb_i_reset[673]                      =   1'b0;
assign   tb_i_sop[673]                        =   1'b0;
assign   tb_i_key_update[673]                 =   1'b0;
assign   tb_i_key[673]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[673]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[673]               =   1'b0;
assign   tb_i_rf_static_encrypt[673]          =   1'b1;
assign   tb_i_clear_fault_flags[673]          =   1'b0;
assign   tb_i_rf_static_aad_length[673]       =   64'h0000000000000100;
assign   tb_i_aad[673]                        =   tb_i_aad[672];
assign   tb_i_rf_static_plaintext_length[673] =   64'h0000000000000280;
assign   tb_i_plaintext[673]                  =   tb_i_plaintext[672];
assign   tb_o_valid[673]                      =   1'b0;
assign   tb_o_sop[673]                        =   1'b0;
assign   tb_o_ciphertext[673]                 =   tb_o_ciphertext[672];
assign   tb_o_tag_ready[673]                  =   1'b0;
assign   tb_o_tag[673]                        =   tb_o_tag[672];

// CLK no. 674/1240
// *************************************************
assign   tb_i_valid[674]                      =   1'b0;
assign   tb_i_reset[674]                      =   1'b0;
assign   tb_i_sop[674]                        =   1'b0;
assign   tb_i_key_update[674]                 =   1'b0;
assign   tb_i_key[674]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[674]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[674]               =   1'b0;
assign   tb_i_rf_static_encrypt[674]          =   1'b1;
assign   tb_i_clear_fault_flags[674]          =   1'b0;
assign   tb_i_rf_static_aad_length[674]       =   64'h0000000000000100;
assign   tb_i_aad[674]                        =   tb_i_aad[673];
assign   tb_i_rf_static_plaintext_length[674] =   64'h0000000000000280;
assign   tb_i_plaintext[674]                  =   tb_i_plaintext[673];
assign   tb_o_valid[674]                      =   1'b0;
assign   tb_o_sop[674]                        =   1'b0;
assign   tb_o_ciphertext[674]                 =   tb_o_ciphertext[673];
assign   tb_o_tag_ready[674]                  =   1'b0;
assign   tb_o_tag[674]                        =   tb_o_tag[673];

// CLK no. 675/1240
// *************************************************
assign   tb_i_valid[675]                      =   1'b0;
assign   tb_i_reset[675]                      =   1'b0;
assign   tb_i_sop[675]                        =   1'b0;
assign   tb_i_key_update[675]                 =   1'b0;
assign   tb_i_key[675]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[675]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[675]               =   1'b0;
assign   tb_i_rf_static_encrypt[675]          =   1'b1;
assign   tb_i_clear_fault_flags[675]          =   1'b0;
assign   tb_i_rf_static_aad_length[675]       =   64'h0000000000000100;
assign   tb_i_aad[675]                        =   tb_i_aad[674];
assign   tb_i_rf_static_plaintext_length[675] =   64'h0000000000000280;
assign   tb_i_plaintext[675]                  =   tb_i_plaintext[674];
assign   tb_o_valid[675]                      =   1'b0;
assign   tb_o_sop[675]                        =   1'b0;
assign   tb_o_ciphertext[675]                 =   tb_o_ciphertext[674];
assign   tb_o_tag_ready[675]                  =   1'b0;
assign   tb_o_tag[675]                        =   tb_o_tag[674];

// CLK no. 676/1240
// *************************************************
assign   tb_i_valid[676]                      =   1'b0;
assign   tb_i_reset[676]                      =   1'b0;
assign   tb_i_sop[676]                        =   1'b0;
assign   tb_i_key_update[676]                 =   1'b0;
assign   tb_i_key[676]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[676]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[676]               =   1'b0;
assign   tb_i_rf_static_encrypt[676]          =   1'b1;
assign   tb_i_clear_fault_flags[676]          =   1'b0;
assign   tb_i_rf_static_aad_length[676]       =   64'h0000000000000100;
assign   tb_i_aad[676]                        =   tb_i_aad[675];
assign   tb_i_rf_static_plaintext_length[676] =   64'h0000000000000280;
assign   tb_i_plaintext[676]                  =   tb_i_plaintext[675];
assign   tb_o_valid[676]                      =   1'b0;
assign   tb_o_sop[676]                        =   1'b0;
assign   tb_o_ciphertext[676]                 =   tb_o_ciphertext[675];
assign   tb_o_tag_ready[676]                  =   1'b0;
assign   tb_o_tag[676]                        =   tb_o_tag[675];

// CLK no. 677/1240
// *************************************************
assign   tb_i_valid[677]                      =   1'b0;
assign   tb_i_reset[677]                      =   1'b0;
assign   tb_i_sop[677]                        =   1'b0;
assign   tb_i_key_update[677]                 =   1'b0;
assign   tb_i_key[677]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[677]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[677]               =   1'b0;
assign   tb_i_rf_static_encrypt[677]          =   1'b1;
assign   tb_i_clear_fault_flags[677]          =   1'b0;
assign   tb_i_rf_static_aad_length[677]       =   64'h0000000000000100;
assign   tb_i_aad[677]                        =   tb_i_aad[676];
assign   tb_i_rf_static_plaintext_length[677] =   64'h0000000000000280;
assign   tb_i_plaintext[677]                  =   tb_i_plaintext[676];
assign   tb_o_valid[677]                      =   1'b0;
assign   tb_o_sop[677]                        =   1'b0;
assign   tb_o_ciphertext[677]                 =   tb_o_ciphertext[676];
assign   tb_o_tag_ready[677]                  =   1'b0;
assign   tb_o_tag[677]                        =   tb_o_tag[676];

// CLK no. 678/1240
// *************************************************
assign   tb_i_valid[678]                      =   1'b0;
assign   tb_i_reset[678]                      =   1'b0;
assign   tb_i_sop[678]                        =   1'b0;
assign   tb_i_key_update[678]                 =   1'b0;
assign   tb_i_key[678]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[678]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[678]               =   1'b0;
assign   tb_i_rf_static_encrypt[678]          =   1'b1;
assign   tb_i_clear_fault_flags[678]          =   1'b0;
assign   tb_i_rf_static_aad_length[678]       =   64'h0000000000000100;
assign   tb_i_aad[678]                        =   tb_i_aad[677];
assign   tb_i_rf_static_plaintext_length[678] =   64'h0000000000000280;
assign   tb_i_plaintext[678]                  =   tb_i_plaintext[677];
assign   tb_o_valid[678]                      =   1'b0;
assign   tb_o_sop[678]                        =   1'b0;
assign   tb_o_ciphertext[678]                 =   tb_o_ciphertext[677];
assign   tb_o_tag_ready[678]                  =   1'b0;
assign   tb_o_tag[678]                        =   tb_o_tag[677];

// CLK no. 679/1240
// *************************************************
assign   tb_i_valid[679]                      =   1'b0;
assign   tb_i_reset[679]                      =   1'b0;
assign   tb_i_sop[679]                        =   1'b0;
assign   tb_i_key_update[679]                 =   1'b0;
assign   tb_i_key[679]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[679]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[679]               =   1'b0;
assign   tb_i_rf_static_encrypt[679]          =   1'b1;
assign   tb_i_clear_fault_flags[679]          =   1'b0;
assign   tb_i_rf_static_aad_length[679]       =   64'h0000000000000100;
assign   tb_i_aad[679]                        =   tb_i_aad[678];
assign   tb_i_rf_static_plaintext_length[679] =   64'h0000000000000280;
assign   tb_i_plaintext[679]                  =   tb_i_plaintext[678];
assign   tb_o_valid[679]                      =   1'b0;
assign   tb_o_sop[679]                        =   1'b0;
assign   tb_o_ciphertext[679]                 =   tb_o_ciphertext[678];
assign   tb_o_tag_ready[679]                  =   1'b0;
assign   tb_o_tag[679]                        =   tb_o_tag[678];

// CLK no. 680/1240
// *************************************************
assign   tb_i_valid[680]                      =   1'b0;
assign   tb_i_reset[680]                      =   1'b0;
assign   tb_i_sop[680]                        =   1'b0;
assign   tb_i_key_update[680]                 =   1'b0;
assign   tb_i_key[680]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[680]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[680]               =   1'b0;
assign   tb_i_rf_static_encrypt[680]          =   1'b1;
assign   tb_i_clear_fault_flags[680]          =   1'b0;
assign   tb_i_rf_static_aad_length[680]       =   64'h0000000000000100;
assign   tb_i_aad[680]                        =   tb_i_aad[679];
assign   tb_i_rf_static_plaintext_length[680] =   64'h0000000000000280;
assign   tb_i_plaintext[680]                  =   tb_i_plaintext[679];
assign   tb_o_valid[680]                      =   1'b0;
assign   tb_o_sop[680]                        =   1'b0;
assign   tb_o_ciphertext[680]                 =   tb_o_ciphertext[679];
assign   tb_o_tag_ready[680]                  =   1'b0;
assign   tb_o_tag[680]                        =   tb_o_tag[679];

// CLK no. 681/1240
// *************************************************
assign   tb_i_valid[681]                      =   1'b0;
assign   tb_i_reset[681]                      =   1'b0;
assign   tb_i_sop[681]                        =   1'b0;
assign   tb_i_key_update[681]                 =   1'b0;
assign   tb_i_key[681]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[681]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[681]               =   1'b0;
assign   tb_i_rf_static_encrypt[681]          =   1'b1;
assign   tb_i_clear_fault_flags[681]          =   1'b0;
assign   tb_i_rf_static_aad_length[681]       =   64'h0000000000000100;
assign   tb_i_aad[681]                        =   tb_i_aad[680];
assign   tb_i_rf_static_plaintext_length[681] =   64'h0000000000000280;
assign   tb_i_plaintext[681]                  =   tb_i_plaintext[680];
assign   tb_o_valid[681]                      =   1'b0;
assign   tb_o_sop[681]                        =   1'b0;
assign   tb_o_ciphertext[681]                 =   tb_o_ciphertext[680];
assign   tb_o_tag_ready[681]                  =   1'b0;
assign   tb_o_tag[681]                        =   tb_o_tag[680];

// CLK no. 682/1240
// *************************************************
assign   tb_i_valid[682]                      =   1'b0;
assign   tb_i_reset[682]                      =   1'b0;
assign   tb_i_sop[682]                        =   1'b0;
assign   tb_i_key_update[682]                 =   1'b0;
assign   tb_i_key[682]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[682]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[682]               =   1'b0;
assign   tb_i_rf_static_encrypt[682]          =   1'b1;
assign   tb_i_clear_fault_flags[682]          =   1'b0;
assign   tb_i_rf_static_aad_length[682]       =   64'h0000000000000100;
assign   tb_i_aad[682]                        =   tb_i_aad[681];
assign   tb_i_rf_static_plaintext_length[682] =   64'h0000000000000280;
assign   tb_i_plaintext[682]                  =   tb_i_plaintext[681];
assign   tb_o_valid[682]                      =   1'b0;
assign   tb_o_sop[682]                        =   1'b0;
assign   tb_o_ciphertext[682]                 =   tb_o_ciphertext[681];
assign   tb_o_tag_ready[682]                  =   1'b0;
assign   tb_o_tag[682]                        =   tb_o_tag[681];

// CLK no. 683/1240
// *************************************************
assign   tb_i_valid[683]                      =   1'b0;
assign   tb_i_reset[683]                      =   1'b0;
assign   tb_i_sop[683]                        =   1'b0;
assign   tb_i_key_update[683]                 =   1'b0;
assign   tb_i_key[683]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[683]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[683]               =   1'b0;
assign   tb_i_rf_static_encrypt[683]          =   1'b1;
assign   tb_i_clear_fault_flags[683]          =   1'b0;
assign   tb_i_rf_static_aad_length[683]       =   64'h0000000000000100;
assign   tb_i_aad[683]                        =   tb_i_aad[682];
assign   tb_i_rf_static_plaintext_length[683] =   64'h0000000000000280;
assign   tb_i_plaintext[683]                  =   tb_i_plaintext[682];
assign   tb_o_valid[683]                      =   1'b0;
assign   tb_o_sop[683]                        =   1'b0;
assign   tb_o_ciphertext[683]                 =   tb_o_ciphertext[682];
assign   tb_o_tag_ready[683]                  =   1'b0;
assign   tb_o_tag[683]                        =   tb_o_tag[682];

// CLK no. 684/1240
// *************************************************
assign   tb_i_valid[684]                      =   1'b0;
assign   tb_i_reset[684]                      =   1'b0;
assign   tb_i_sop[684]                        =   1'b0;
assign   tb_i_key_update[684]                 =   1'b0;
assign   tb_i_key[684]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[684]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[684]               =   1'b0;
assign   tb_i_rf_static_encrypt[684]          =   1'b1;
assign   tb_i_clear_fault_flags[684]          =   1'b0;
assign   tb_i_rf_static_aad_length[684]       =   64'h0000000000000100;
assign   tb_i_aad[684]                        =   tb_i_aad[683];
assign   tb_i_rf_static_plaintext_length[684] =   64'h0000000000000280;
assign   tb_i_plaintext[684]                  =   tb_i_plaintext[683];
assign   tb_o_valid[684]                      =   1'b0;
assign   tb_o_sop[684]                        =   1'b0;
assign   tb_o_ciphertext[684]                 =   tb_o_ciphertext[683];
assign   tb_o_tag_ready[684]                  =   1'b0;
assign   tb_o_tag[684]                        =   tb_o_tag[683];

// CLK no. 685/1240
// *************************************************
assign   tb_i_valid[685]                      =   1'b0;
assign   tb_i_reset[685]                      =   1'b0;
assign   tb_i_sop[685]                        =   1'b0;
assign   tb_i_key_update[685]                 =   1'b0;
assign   tb_i_key[685]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[685]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[685]               =   1'b0;
assign   tb_i_rf_static_encrypt[685]          =   1'b1;
assign   tb_i_clear_fault_flags[685]          =   1'b0;
assign   tb_i_rf_static_aad_length[685]       =   64'h0000000000000100;
assign   tb_i_aad[685]                        =   tb_i_aad[684];
assign   tb_i_rf_static_plaintext_length[685] =   64'h0000000000000280;
assign   tb_i_plaintext[685]                  =   tb_i_plaintext[684];
assign   tb_o_valid[685]                      =   1'b0;
assign   tb_o_sop[685]                        =   1'b0;
assign   tb_o_ciphertext[685]                 =   tb_o_ciphertext[684];
assign   tb_o_tag_ready[685]                  =   1'b0;
assign   tb_o_tag[685]                        =   tb_o_tag[684];

// CLK no. 686/1240
// *************************************************
assign   tb_i_valid[686]                      =   1'b0;
assign   tb_i_reset[686]                      =   1'b0;
assign   tb_i_sop[686]                        =   1'b0;
assign   tb_i_key_update[686]                 =   1'b0;
assign   tb_i_key[686]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[686]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[686]               =   1'b0;
assign   tb_i_rf_static_encrypt[686]          =   1'b1;
assign   tb_i_clear_fault_flags[686]          =   1'b0;
assign   tb_i_rf_static_aad_length[686]       =   64'h0000000000000100;
assign   tb_i_aad[686]                        =   tb_i_aad[685];
assign   tb_i_rf_static_plaintext_length[686] =   64'h0000000000000280;
assign   tb_i_plaintext[686]                  =   tb_i_plaintext[685];
assign   tb_o_valid[686]                      =   1'b0;
assign   tb_o_sop[686]                        =   1'b0;
assign   tb_o_ciphertext[686]                 =   tb_o_ciphertext[685];
assign   tb_o_tag_ready[686]                  =   1'b0;
assign   tb_o_tag[686]                        =   tb_o_tag[685];

// CLK no. 687/1240
// *************************************************
assign   tb_i_valid[687]                      =   1'b0;
assign   tb_i_reset[687]                      =   1'b0;
assign   tb_i_sop[687]                        =   1'b0;
assign   tb_i_key_update[687]                 =   1'b0;
assign   tb_i_key[687]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[687]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[687]               =   1'b0;
assign   tb_i_rf_static_encrypt[687]          =   1'b1;
assign   tb_i_clear_fault_flags[687]          =   1'b0;
assign   tb_i_rf_static_aad_length[687]       =   64'h0000000000000100;
assign   tb_i_aad[687]                        =   tb_i_aad[686];
assign   tb_i_rf_static_plaintext_length[687] =   64'h0000000000000280;
assign   tb_i_plaintext[687]                  =   tb_i_plaintext[686];
assign   tb_o_valid[687]                      =   1'b0;
assign   tb_o_sop[687]                        =   1'b0;
assign   tb_o_ciphertext[687]                 =   tb_o_ciphertext[686];
assign   tb_o_tag_ready[687]                  =   1'b0;
assign   tb_o_tag[687]                        =   tb_o_tag[686];

// CLK no. 688/1240
// *************************************************
assign   tb_i_valid[688]                      =   1'b0;
assign   tb_i_reset[688]                      =   1'b0;
assign   tb_i_sop[688]                        =   1'b0;
assign   tb_i_key_update[688]                 =   1'b0;
assign   tb_i_key[688]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[688]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[688]               =   1'b0;
assign   tb_i_rf_static_encrypt[688]          =   1'b1;
assign   tb_i_clear_fault_flags[688]          =   1'b0;
assign   tb_i_rf_static_aad_length[688]       =   64'h0000000000000100;
assign   tb_i_aad[688]                        =   tb_i_aad[687];
assign   tb_i_rf_static_plaintext_length[688] =   64'h0000000000000280;
assign   tb_i_plaintext[688]                  =   tb_i_plaintext[687];
assign   tb_o_valid[688]                      =   1'b0;
assign   tb_o_sop[688]                        =   1'b0;
assign   tb_o_ciphertext[688]                 =   tb_o_ciphertext[687];
assign   tb_o_tag_ready[688]                  =   1'b0;
assign   tb_o_tag[688]                        =   tb_o_tag[687];

// CLK no. 689/1240
// *************************************************
assign   tb_i_valid[689]                      =   1'b0;
assign   tb_i_reset[689]                      =   1'b0;
assign   tb_i_sop[689]                        =   1'b0;
assign   tb_i_key_update[689]                 =   1'b0;
assign   tb_i_key[689]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[689]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[689]               =   1'b0;
assign   tb_i_rf_static_encrypt[689]          =   1'b1;
assign   tb_i_clear_fault_flags[689]          =   1'b0;
assign   tb_i_rf_static_aad_length[689]       =   64'h0000000000000100;
assign   tb_i_aad[689]                        =   tb_i_aad[688];
assign   tb_i_rf_static_plaintext_length[689] =   64'h0000000000000280;
assign   tb_i_plaintext[689]                  =   tb_i_plaintext[688];
assign   tb_o_valid[689]                      =   1'b0;
assign   tb_o_sop[689]                        =   1'b0;
assign   tb_o_ciphertext[689]                 =   tb_o_ciphertext[688];
assign   tb_o_tag_ready[689]                  =   1'b0;
assign   tb_o_tag[689]                        =   tb_o_tag[688];

// CLK no. 690/1240
// *************************************************
assign   tb_i_valid[690]                      =   1'b0;
assign   tb_i_reset[690]                      =   1'b0;
assign   tb_i_sop[690]                        =   1'b0;
assign   tb_i_key_update[690]                 =   1'b0;
assign   tb_i_key[690]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[690]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[690]               =   1'b0;
assign   tb_i_rf_static_encrypt[690]          =   1'b1;
assign   tb_i_clear_fault_flags[690]          =   1'b0;
assign   tb_i_rf_static_aad_length[690]       =   64'h0000000000000100;
assign   tb_i_aad[690]                        =   tb_i_aad[689];
assign   tb_i_rf_static_plaintext_length[690] =   64'h0000000000000280;
assign   tb_i_plaintext[690]                  =   tb_i_plaintext[689];
assign   tb_o_valid[690]                      =   1'b0;
assign   tb_o_sop[690]                        =   1'b0;
assign   tb_o_ciphertext[690]                 =   tb_o_ciphertext[689];
assign   tb_o_tag_ready[690]                  =   1'b0;
assign   tb_o_tag[690]                        =   tb_o_tag[689];

// CLK no. 691/1240
// *************************************************
assign   tb_i_valid[691]                      =   1'b0;
assign   tb_i_reset[691]                      =   1'b0;
assign   tb_i_sop[691]                        =   1'b0;
assign   tb_i_key_update[691]                 =   1'b0;
assign   tb_i_key[691]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[691]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[691]               =   1'b0;
assign   tb_i_rf_static_encrypt[691]          =   1'b1;
assign   tb_i_clear_fault_flags[691]          =   1'b0;
assign   tb_i_rf_static_aad_length[691]       =   64'h0000000000000100;
assign   tb_i_aad[691]                        =   tb_i_aad[690];
assign   tb_i_rf_static_plaintext_length[691] =   64'h0000000000000280;
assign   tb_i_plaintext[691]                  =   tb_i_plaintext[690];
assign   tb_o_valid[691]                      =   1'b0;
assign   tb_o_sop[691]                        =   1'b0;
assign   tb_o_ciphertext[691]                 =   tb_o_ciphertext[690];
assign   tb_o_tag_ready[691]                  =   1'b0;
assign   tb_o_tag[691]                        =   tb_o_tag[690];

// CLK no. 692/1240
// *************************************************
assign   tb_i_valid[692]                      =   1'b0;
assign   tb_i_reset[692]                      =   1'b0;
assign   tb_i_sop[692]                        =   1'b0;
assign   tb_i_key_update[692]                 =   1'b0;
assign   tb_i_key[692]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[692]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[692]               =   1'b0;
assign   tb_i_rf_static_encrypt[692]          =   1'b1;
assign   tb_i_clear_fault_flags[692]          =   1'b0;
assign   tb_i_rf_static_aad_length[692]       =   64'h0000000000000100;
assign   tb_i_aad[692]                        =   tb_i_aad[691];
assign   tb_i_rf_static_plaintext_length[692] =   64'h0000000000000280;
assign   tb_i_plaintext[692]                  =   tb_i_plaintext[691];
assign   tb_o_valid[692]                      =   1'b0;
assign   tb_o_sop[692]                        =   1'b0;
assign   tb_o_ciphertext[692]                 =   tb_o_ciphertext[691];
assign   tb_o_tag_ready[692]                  =   1'b0;
assign   tb_o_tag[692]                        =   tb_o_tag[691];

// CLK no. 693/1240
// *************************************************
assign   tb_i_valid[693]                      =   1'b0;
assign   tb_i_reset[693]                      =   1'b0;
assign   tb_i_sop[693]                        =   1'b0;
assign   tb_i_key_update[693]                 =   1'b0;
assign   tb_i_key[693]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[693]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[693]               =   1'b0;
assign   tb_i_rf_static_encrypt[693]          =   1'b1;
assign   tb_i_clear_fault_flags[693]          =   1'b0;
assign   tb_i_rf_static_aad_length[693]       =   64'h0000000000000100;
assign   tb_i_aad[693]                        =   tb_i_aad[692];
assign   tb_i_rf_static_plaintext_length[693] =   64'h0000000000000280;
assign   tb_i_plaintext[693]                  =   tb_i_plaintext[692];
assign   tb_o_valid[693]                      =   1'b0;
assign   tb_o_sop[693]                        =   1'b0;
assign   tb_o_ciphertext[693]                 =   tb_o_ciphertext[692];
assign   tb_o_tag_ready[693]                  =   1'b0;
assign   tb_o_tag[693]                        =   tb_o_tag[692];

// CLK no. 694/1240
// *************************************************
assign   tb_i_valid[694]                      =   1'b0;
assign   tb_i_reset[694]                      =   1'b0;
assign   tb_i_sop[694]                        =   1'b0;
assign   tb_i_key_update[694]                 =   1'b0;
assign   tb_i_key[694]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[694]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[694]               =   1'b0;
assign   tb_i_rf_static_encrypt[694]          =   1'b1;
assign   tb_i_clear_fault_flags[694]          =   1'b0;
assign   tb_i_rf_static_aad_length[694]       =   64'h0000000000000100;
assign   tb_i_aad[694]                        =   tb_i_aad[693];
assign   tb_i_rf_static_plaintext_length[694] =   64'h0000000000000280;
assign   tb_i_plaintext[694]                  =   tb_i_plaintext[693];
assign   tb_o_valid[694]                      =   1'b0;
assign   tb_o_sop[694]                        =   1'b0;
assign   tb_o_ciphertext[694]                 =   tb_o_ciphertext[693];
assign   tb_o_tag_ready[694]                  =   1'b0;
assign   tb_o_tag[694]                        =   tb_o_tag[693];

// CLK no. 695/1240
// *************************************************
assign   tb_i_valid[695]                      =   1'b0;
assign   tb_i_reset[695]                      =   1'b0;
assign   tb_i_sop[695]                        =   1'b0;
assign   tb_i_key_update[695]                 =   1'b0;
assign   tb_i_key[695]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[695]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[695]               =   1'b0;
assign   tb_i_rf_static_encrypt[695]          =   1'b1;
assign   tb_i_clear_fault_flags[695]          =   1'b0;
assign   tb_i_rf_static_aad_length[695]       =   64'h0000000000000100;
assign   tb_i_aad[695]                        =   tb_i_aad[694];
assign   tb_i_rf_static_plaintext_length[695] =   64'h0000000000000280;
assign   tb_i_plaintext[695]                  =   tb_i_plaintext[694];
assign   tb_o_valid[695]                      =   1'b0;
assign   tb_o_sop[695]                        =   1'b0;
assign   tb_o_ciphertext[695]                 =   tb_o_ciphertext[694];
assign   tb_o_tag_ready[695]                  =   1'b0;
assign   tb_o_tag[695]                        =   tb_o_tag[694];

// CLK no. 696/1240
// *************************************************
assign   tb_i_valid[696]                      =   1'b0;
assign   tb_i_reset[696]                      =   1'b0;
assign   tb_i_sop[696]                        =   1'b0;
assign   tb_i_key_update[696]                 =   1'b0;
assign   tb_i_key[696]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[696]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[696]               =   1'b0;
assign   tb_i_rf_static_encrypt[696]          =   1'b1;
assign   tb_i_clear_fault_flags[696]          =   1'b0;
assign   tb_i_rf_static_aad_length[696]       =   64'h0000000000000100;
assign   tb_i_aad[696]                        =   tb_i_aad[695];
assign   tb_i_rf_static_plaintext_length[696] =   64'h0000000000000280;
assign   tb_i_plaintext[696]                  =   tb_i_plaintext[695];
assign   tb_o_valid[696]                      =   1'b1;
assign   tb_o_sop[696]                        =   1'b1;
assign   tb_o_ciphertext[696]                 =   256'h5f6c8874c6372f94a736abfe8e18b2d461f7eaafff6111cfd642bd36c6ee4b3d;
assign   tb_o_tag_ready[696]                  =   1'b0;
assign   tb_o_tag[696]                        =   tb_o_tag[695];

// CLK no. 697/1240
// *************************************************
assign   tb_i_valid[697]                      =   1'b0;
assign   tb_i_reset[697]                      =   1'b0;
assign   tb_i_sop[697]                        =   1'b0;
assign   tb_i_key_update[697]                 =   1'b0;
assign   tb_i_key[697]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[697]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[697]               =   1'b0;
assign   tb_i_rf_static_encrypt[697]          =   1'b1;
assign   tb_i_clear_fault_flags[697]          =   1'b0;
assign   tb_i_rf_static_aad_length[697]       =   64'h0000000000000100;
assign   tb_i_aad[697]                        =   tb_i_aad[696];
assign   tb_i_rf_static_plaintext_length[697] =   64'h0000000000000280;
assign   tb_i_plaintext[697]                  =   tb_i_plaintext[696];
assign   tb_o_valid[697]                      =   1'b1;
assign   tb_o_sop[697]                        =   1'b0;
assign   tb_o_ciphertext[697]                 =   256'h8927a6fa5395e491b03622e6b6ce0846dc5b73929c20a9abc78cc9c3dddae01e;
assign   tb_o_tag_ready[697]                  =   1'b0;
assign   tb_o_tag[697]                        =   tb_o_tag[696];

// CLK no. 698/1240
// *************************************************
assign   tb_i_valid[698]                      =   1'b0;
assign   tb_i_reset[698]                      =   1'b0;
assign   tb_i_sop[698]                        =   1'b0;
assign   tb_i_key_update[698]                 =   1'b0;
assign   tb_i_key[698]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[698]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[698]               =   1'b0;
assign   tb_i_rf_static_encrypt[698]          =   1'b1;
assign   tb_i_clear_fault_flags[698]          =   1'b0;
assign   tb_i_rf_static_aad_length[698]       =   64'h0000000000000100;
assign   tb_i_aad[698]                        =   tb_i_aad[697];
assign   tb_i_rf_static_plaintext_length[698] =   64'h0000000000000280;
assign   tb_i_plaintext[698]                  =   tb_i_plaintext[697];
assign   tb_o_valid[698]                      =   1'b1;
assign   tb_o_sop[698]                        =   1'b0;
assign   tb_o_ciphertext[698]                 =   256'hbbce0932f5d92899d53305dc3bafa1f8;
assign   tb_o_tag_ready[698]                  =   1'b0;
assign   tb_o_tag[698]                        =   tb_o_tag[697];

// CLK no. 699/1240
// *************************************************
assign   tb_i_valid[699]                      =   1'b0;
assign   tb_i_reset[699]                      =   1'b0;
assign   tb_i_sop[699]                        =   1'b0;
assign   tb_i_key_update[699]                 =   1'b0;
assign   tb_i_key[699]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[699]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[699]               =   1'b0;
assign   tb_i_rf_static_encrypt[699]          =   1'b1;
assign   tb_i_clear_fault_flags[699]          =   1'b0;
assign   tb_i_rf_static_aad_length[699]       =   64'h0000000000000100;
assign   tb_i_aad[699]                        =   tb_i_aad[698];
assign   tb_i_rf_static_plaintext_length[699] =   64'h0000000000000280;
assign   tb_i_plaintext[699]                  =   tb_i_plaintext[698];
assign   tb_o_valid[699]                      =   1'b0;
assign   tb_o_sop[699]                        =   1'b0;
assign   tb_o_ciphertext[699]                 =   tb_o_ciphertext[698];
assign   tb_o_tag_ready[699]                  =   1'b0;
assign   tb_o_tag[699]                        =   tb_o_tag[698];

// CLK no. 700/1240
// *************************************************
assign   tb_i_valid[700]                      =   1'b0;
assign   tb_i_reset[700]                      =   1'b0;
assign   tb_i_sop[700]                        =   1'b0;
assign   tb_i_key_update[700]                 =   1'b0;
assign   tb_i_key[700]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[700]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[700]               =   1'b0;
assign   tb_i_rf_static_encrypt[700]          =   1'b1;
assign   tb_i_clear_fault_flags[700]          =   1'b0;
assign   tb_i_rf_static_aad_length[700]       =   64'h0000000000000100;
assign   tb_i_aad[700]                        =   tb_i_aad[699];
assign   tb_i_rf_static_plaintext_length[700] =   64'h0000000000000280;
assign   tb_i_plaintext[700]                  =   tb_i_plaintext[699];
assign   tb_o_valid[700]                      =   1'b0;
assign   tb_o_sop[700]                        =   1'b0;
assign   tb_o_ciphertext[700]                 =   tb_o_ciphertext[699];
assign   tb_o_tag_ready[700]                  =   1'b0;
assign   tb_o_tag[700]                        =   tb_o_tag[699];

// CLK no. 701/1240
// *************************************************
assign   tb_i_valid[701]                      =   1'b0;
assign   tb_i_reset[701]                      =   1'b0;
assign   tb_i_sop[701]                        =   1'b0;
assign   tb_i_key_update[701]                 =   1'b0;
assign   tb_i_key[701]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[701]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[701]               =   1'b0;
assign   tb_i_rf_static_encrypt[701]          =   1'b1;
assign   tb_i_clear_fault_flags[701]          =   1'b0;
assign   tb_i_rf_static_aad_length[701]       =   64'h0000000000000100;
assign   tb_i_aad[701]                        =   tb_i_aad[700];
assign   tb_i_rf_static_plaintext_length[701] =   64'h0000000000000280;
assign   tb_i_plaintext[701]                  =   tb_i_plaintext[700];
assign   tb_o_valid[701]                      =   1'b0;
assign   tb_o_sop[701]                        =   1'b0;
assign   tb_o_ciphertext[701]                 =   tb_o_ciphertext[700];
assign   tb_o_tag_ready[701]                  =   1'b0;
assign   tb_o_tag[701]                        =   tb_o_tag[700];

// CLK no. 702/1240
// *************************************************
assign   tb_i_valid[702]                      =   1'b0;
assign   tb_i_reset[702]                      =   1'b0;
assign   tb_i_sop[702]                        =   1'b0;
assign   tb_i_key_update[702]                 =   1'b0;
assign   tb_i_key[702]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[702]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[702]               =   1'b0;
assign   tb_i_rf_static_encrypt[702]          =   1'b1;
assign   tb_i_clear_fault_flags[702]          =   1'b0;
assign   tb_i_rf_static_aad_length[702]       =   64'h0000000000000100;
assign   tb_i_aad[702]                        =   tb_i_aad[701];
assign   tb_i_rf_static_plaintext_length[702] =   64'h0000000000000280;
assign   tb_i_plaintext[702]                  =   tb_i_plaintext[701];
assign   tb_o_valid[702]                      =   1'b0;
assign   tb_o_sop[702]                        =   1'b0;
assign   tb_o_ciphertext[702]                 =   tb_o_ciphertext[701];
assign   tb_o_tag_ready[702]                  =   1'b0;
assign   tb_o_tag[702]                        =   tb_o_tag[701];

// CLK no. 703/1240
// *************************************************
assign   tb_i_valid[703]                      =   1'b0;
assign   tb_i_reset[703]                      =   1'b0;
assign   tb_i_sop[703]                        =   1'b0;
assign   tb_i_key_update[703]                 =   1'b0;
assign   tb_i_key[703]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[703]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[703]               =   1'b0;
assign   tb_i_rf_static_encrypt[703]          =   1'b1;
assign   tb_i_clear_fault_flags[703]          =   1'b0;
assign   tb_i_rf_static_aad_length[703]       =   64'h0000000000000100;
assign   tb_i_aad[703]                        =   tb_i_aad[702];
assign   tb_i_rf_static_plaintext_length[703] =   64'h0000000000000280;
assign   tb_i_plaintext[703]                  =   tb_i_plaintext[702];
assign   tb_o_valid[703]                      =   1'b0;
assign   tb_o_sop[703]                        =   1'b0;
assign   tb_o_ciphertext[703]                 =   tb_o_ciphertext[702];
assign   tb_o_tag_ready[703]                  =   1'b0;
assign   tb_o_tag[703]                        =   tb_o_tag[702];

// CLK no. 704/1240
// *************************************************
assign   tb_i_valid[704]                      =   1'b0;
assign   tb_i_reset[704]                      =   1'b0;
assign   tb_i_sop[704]                        =   1'b0;
assign   tb_i_key_update[704]                 =   1'b0;
assign   tb_i_key[704]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[704]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[704]               =   1'b0;
assign   tb_i_rf_static_encrypt[704]          =   1'b1;
assign   tb_i_clear_fault_flags[704]          =   1'b0;
assign   tb_i_rf_static_aad_length[704]       =   64'h0000000000000100;
assign   tb_i_aad[704]                        =   tb_i_aad[703];
assign   tb_i_rf_static_plaintext_length[704] =   64'h0000000000000280;
assign   tb_i_plaintext[704]                  =   tb_i_plaintext[703];
assign   tb_o_valid[704]                      =   1'b0;
assign   tb_o_sop[704]                        =   1'b0;
assign   tb_o_ciphertext[704]                 =   tb_o_ciphertext[703];
assign   tb_o_tag_ready[704]                  =   1'b0;
assign   tb_o_tag[704]                        =   tb_o_tag[703];

// CLK no. 705/1240
// *************************************************
assign   tb_i_valid[705]                      =   1'b0;
assign   tb_i_reset[705]                      =   1'b0;
assign   tb_i_sop[705]                        =   1'b0;
assign   tb_i_key_update[705]                 =   1'b0;
assign   tb_i_key[705]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[705]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[705]               =   1'b0;
assign   tb_i_rf_static_encrypt[705]          =   1'b1;
assign   tb_i_clear_fault_flags[705]          =   1'b0;
assign   tb_i_rf_static_aad_length[705]       =   64'h0000000000000100;
assign   tb_i_aad[705]                        =   tb_i_aad[704];
assign   tb_i_rf_static_plaintext_length[705] =   64'h0000000000000280;
assign   tb_i_plaintext[705]                  =   tb_i_plaintext[704];
assign   tb_o_valid[705]                      =   1'b0;
assign   tb_o_sop[705]                        =   1'b0;
assign   tb_o_ciphertext[705]                 =   tb_o_ciphertext[704];
assign   tb_o_tag_ready[705]                  =   1'b0;
assign   tb_o_tag[705]                        =   tb_o_tag[704];

// CLK no. 706/1240
// *************************************************
assign   tb_i_valid[706]                      =   1'b0;
assign   tb_i_reset[706]                      =   1'b0;
assign   tb_i_sop[706]                        =   1'b0;
assign   tb_i_key_update[706]                 =   1'b0;
assign   tb_i_key[706]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[706]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[706]               =   1'b0;
assign   tb_i_rf_static_encrypt[706]          =   1'b1;
assign   tb_i_clear_fault_flags[706]          =   1'b0;
assign   tb_i_rf_static_aad_length[706]       =   64'h0000000000000100;
assign   tb_i_aad[706]                        =   tb_i_aad[705];
assign   tb_i_rf_static_plaintext_length[706] =   64'h0000000000000280;
assign   tb_i_plaintext[706]                  =   tb_i_plaintext[705];
assign   tb_o_valid[706]                      =   1'b0;
assign   tb_o_sop[706]                        =   1'b0;
assign   tb_o_ciphertext[706]                 =   tb_o_ciphertext[705];
assign   tb_o_tag_ready[706]                  =   1'b1;
assign   tb_o_tag[706]                        =   128'h55e1e55537e0412315fedf044a8a2cb3;

// CLK no. 707/1240
// *************************************************
assign   tb_i_valid[707]                      =   1'b0;
assign   tb_i_reset[707]                      =   1'b0;
assign   tb_i_sop[707]                        =   1'b0;
assign   tb_i_key_update[707]                 =   1'b0;
assign   tb_i_key[707]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[707]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[707]               =   1'b0;
assign   tb_i_rf_static_encrypt[707]          =   1'b1;
assign   tb_i_clear_fault_flags[707]          =   1'b0;
assign   tb_i_rf_static_aad_length[707]       =   64'h0000000000000100;
assign   tb_i_aad[707]                        =   tb_i_aad[706];
assign   tb_i_rf_static_plaintext_length[707] =   64'h0000000000000280;
assign   tb_i_plaintext[707]                  =   tb_i_plaintext[706];
assign   tb_o_valid[707]                      =   1'b0;
assign   tb_o_sop[707]                        =   1'b0;
assign   tb_o_ciphertext[707]                 =   tb_o_ciphertext[706];
assign   tb_o_tag_ready[707]                  =   1'b0;
assign   tb_o_tag[707]                        =   tb_o_tag[706];

// CLK no. 708/1240
// *************************************************
assign   tb_i_valid[708]                      =   1'b0;
assign   tb_i_reset[708]                      =   1'b0;
assign   tb_i_sop[708]                        =   1'b0;
assign   tb_i_key_update[708]                 =   1'b0;
assign   tb_i_key[708]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[708]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[708]               =   1'b0;
assign   tb_i_rf_static_encrypt[708]          =   1'b1;
assign   tb_i_clear_fault_flags[708]          =   1'b0;
assign   tb_i_rf_static_aad_length[708]       =   64'h0000000000000100;
assign   tb_i_aad[708]                        =   tb_i_aad[707];
assign   tb_i_rf_static_plaintext_length[708] =   64'h0000000000000280;
assign   tb_i_plaintext[708]                  =   tb_i_plaintext[707];
assign   tb_o_valid[708]                      =   1'b0;
assign   tb_o_sop[708]                        =   1'b0;
assign   tb_o_ciphertext[708]                 =   tb_o_ciphertext[707];
assign   tb_o_tag_ready[708]                  =   1'b0;
assign   tb_o_tag[708]                        =   tb_o_tag[707];

// CLK no. 709/1240
// *************************************************
assign   tb_i_valid[709]                      =   1'b0;
assign   tb_i_reset[709]                      =   1'b0;
assign   tb_i_sop[709]                        =   1'b1;
assign   tb_i_key_update[709]                 =   1'b0;
assign   tb_i_key[709]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[709]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[709]               =   1'b0;
assign   tb_i_rf_static_encrypt[709]          =   1'b1;
assign   tb_i_clear_fault_flags[709]          =   1'b0;
assign   tb_i_rf_static_aad_length[709]       =   64'h0000000000000100;
assign   tb_i_aad[709]                        =   tb_i_aad[708];
assign   tb_i_rf_static_plaintext_length[709] =   64'h0000000000000280;
assign   tb_i_plaintext[709]                  =   tb_i_plaintext[708];
assign   tb_o_valid[709]                      =   1'b0;
assign   tb_o_sop[709]                        =   1'b0;
assign   tb_o_ciphertext[709]                 =   tb_o_ciphertext[708];
assign   tb_o_tag_ready[709]                  =   1'b0;
assign   tb_o_tag[709]                        =   tb_o_tag[708];

// CLK no. 710/1240
// *************************************************
assign   tb_i_valid[710]                      =   1'b1;
assign   tb_i_reset[710]                      =   1'b0;
assign   tb_i_sop[710]                        =   1'b0;
assign   tb_i_key_update[710]                 =   1'b0;
assign   tb_i_key[710]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[710]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[710]               =   1'b0;
assign   tb_i_rf_static_encrypt[710]          =   1'b1;
assign   tb_i_clear_fault_flags[710]          =   1'b0;
assign   tb_i_rf_static_aad_length[710]       =   64'h0000000000000100;
assign   tb_i_aad[710]                        =   256'h49791ca2c803fc848efda4b8254219eced351cba9d59cb104c50db294ac1ef3a;
assign   tb_i_rf_static_plaintext_length[710] =   64'h0000000000000280;
assign   tb_i_plaintext[710]                  =   tb_i_plaintext[709];
assign   tb_o_valid[710]                      =   1'b0;
assign   tb_o_sop[710]                        =   1'b0;
assign   tb_o_ciphertext[710]                 =   tb_o_ciphertext[709];
assign   tb_o_tag_ready[710]                  =   1'b0;
assign   tb_o_tag[710]                        =   tb_o_tag[709];

// CLK no. 711/1240
// *************************************************
assign   tb_i_valid[711]                      =   1'b1;
assign   tb_i_reset[711]                      =   1'b0;
assign   tb_i_sop[711]                        =   1'b0;
assign   tb_i_key_update[711]                 =   1'b0;
assign   tb_i_key[711]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[711]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[711]               =   1'b0;
assign   tb_i_rf_static_encrypt[711]          =   1'b1;
assign   tb_i_clear_fault_flags[711]          =   1'b0;
assign   tb_i_rf_static_aad_length[711]       =   64'h0000000000000100;
assign   tb_i_aad[711]                        =   tb_i_aad[710];
assign   tb_i_rf_static_plaintext_length[711] =   64'h0000000000000280;
assign   tb_i_plaintext[711]                  =   256'hc0a37f714106f5b4906704233845dcd18588d17e501e6aa06536f92d29aabdd3;
assign   tb_o_valid[711]                      =   1'b0;
assign   tb_o_sop[711]                        =   1'b0;
assign   tb_o_ciphertext[711]                 =   tb_o_ciphertext[710];
assign   tb_o_tag_ready[711]                  =   1'b0;
assign   tb_o_tag[711]                        =   tb_o_tag[710];

// CLK no. 712/1240
// *************************************************
assign   tb_i_valid[712]                      =   1'b1;
assign   tb_i_reset[712]                      =   1'b0;
assign   tb_i_sop[712]                        =   1'b0;
assign   tb_i_key_update[712]                 =   1'b0;
assign   tb_i_key[712]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[712]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[712]               =   1'b0;
assign   tb_i_rf_static_encrypt[712]          =   1'b1;
assign   tb_i_clear_fault_flags[712]          =   1'b0;
assign   tb_i_rf_static_aad_length[712]       =   64'h0000000000000100;
assign   tb_i_aad[712]                        =   tb_i_aad[711];
assign   tb_i_rf_static_plaintext_length[712] =   64'h0000000000000280;
assign   tb_i_plaintext[712]                  =   256'he082a24d4ede4f18aa319a207a47a0ffbf66cfa274c34cc85e6253b5dd663500;
assign   tb_o_valid[712]                      =   1'b0;
assign   tb_o_sop[712]                        =   1'b0;
assign   tb_o_ciphertext[712]                 =   tb_o_ciphertext[711];
assign   tb_o_tag_ready[712]                  =   1'b0;
assign   tb_o_tag[712]                        =   tb_o_tag[711];

// CLK no. 713/1240
// *************************************************
assign   tb_i_valid[713]                      =   1'b1;
assign   tb_i_reset[713]                      =   1'b0;
assign   tb_i_sop[713]                        =   1'b0;
assign   tb_i_key_update[713]                 =   1'b0;
assign   tb_i_key[713]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[713]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[713]               =   1'b0;
assign   tb_i_rf_static_encrypt[713]          =   1'b1;
assign   tb_i_clear_fault_flags[713]          =   1'b0;
assign   tb_i_rf_static_aad_length[713]       =   64'h0000000000000100;
assign   tb_i_aad[713]                        =   tb_i_aad[712];
assign   tb_i_rf_static_plaintext_length[713] =   64'h0000000000000280;
assign   tb_i_plaintext[713]                  =   256'h2bcaa7c6f891772dcb61d08cfb13f0d8;
assign   tb_o_valid[713]                      =   1'b0;
assign   tb_o_sop[713]                        =   1'b0;
assign   tb_o_ciphertext[713]                 =   tb_o_ciphertext[712];
assign   tb_o_tag_ready[713]                  =   1'b0;
assign   tb_o_tag[713]                        =   tb_o_tag[712];

// CLK no. 714/1240
// *************************************************
assign   tb_i_valid[714]                      =   1'b0;
assign   tb_i_reset[714]                      =   1'b0;
assign   tb_i_sop[714]                        =   1'b0;
assign   tb_i_key_update[714]                 =   1'b0;
assign   tb_i_key[714]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[714]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[714]               =   1'b0;
assign   tb_i_rf_static_encrypt[714]          =   1'b1;
assign   tb_i_clear_fault_flags[714]          =   1'b0;
assign   tb_i_rf_static_aad_length[714]       =   64'h0000000000000100;
assign   tb_i_aad[714]                        =   tb_i_aad[713];
assign   tb_i_rf_static_plaintext_length[714] =   64'h0000000000000280;
assign   tb_i_plaintext[714]                  =   tb_i_plaintext[713];
assign   tb_o_valid[714]                      =   1'b0;
assign   tb_o_sop[714]                        =   1'b0;
assign   tb_o_ciphertext[714]                 =   tb_o_ciphertext[713];
assign   tb_o_tag_ready[714]                  =   1'b0;
assign   tb_o_tag[714]                        =   tb_o_tag[713];

// CLK no. 715/1240
// *************************************************
assign   tb_i_valid[715]                      =   1'b0;
assign   tb_i_reset[715]                      =   1'b0;
assign   tb_i_sop[715]                        =   1'b0;
assign   tb_i_key_update[715]                 =   1'b0;
assign   tb_i_key[715]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[715]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[715]               =   1'b0;
assign   tb_i_rf_static_encrypt[715]          =   1'b1;
assign   tb_i_clear_fault_flags[715]          =   1'b0;
assign   tb_i_rf_static_aad_length[715]       =   64'h0000000000000100;
assign   tb_i_aad[715]                        =   tb_i_aad[714];
assign   tb_i_rf_static_plaintext_length[715] =   64'h0000000000000280;
assign   tb_i_plaintext[715]                  =   tb_i_plaintext[714];
assign   tb_o_valid[715]                      =   1'b0;
assign   tb_o_sop[715]                        =   1'b0;
assign   tb_o_ciphertext[715]                 =   tb_o_ciphertext[714];
assign   tb_o_tag_ready[715]                  =   1'b0;
assign   tb_o_tag[715]                        =   tb_o_tag[714];

// CLK no. 716/1240
// *************************************************
assign   tb_i_valid[716]                      =   1'b0;
assign   tb_i_reset[716]                      =   1'b0;
assign   tb_i_sop[716]                        =   1'b0;
assign   tb_i_key_update[716]                 =   1'b0;
assign   tb_i_key[716]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[716]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[716]               =   1'b0;
assign   tb_i_rf_static_encrypt[716]          =   1'b1;
assign   tb_i_clear_fault_flags[716]          =   1'b0;
assign   tb_i_rf_static_aad_length[716]       =   64'h0000000000000100;
assign   tb_i_aad[716]                        =   tb_i_aad[715];
assign   tb_i_rf_static_plaintext_length[716] =   64'h0000000000000280;
assign   tb_i_plaintext[716]                  =   tb_i_plaintext[715];
assign   tb_o_valid[716]                      =   1'b0;
assign   tb_o_sop[716]                        =   1'b0;
assign   tb_o_ciphertext[716]                 =   tb_o_ciphertext[715];
assign   tb_o_tag_ready[716]                  =   1'b0;
assign   tb_o_tag[716]                        =   tb_o_tag[715];

// CLK no. 717/1240
// *************************************************
assign   tb_i_valid[717]                      =   1'b0;
assign   tb_i_reset[717]                      =   1'b0;
assign   tb_i_sop[717]                        =   1'b0;
assign   tb_i_key_update[717]                 =   1'b0;
assign   tb_i_key[717]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[717]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[717]               =   1'b0;
assign   tb_i_rf_static_encrypt[717]          =   1'b1;
assign   tb_i_clear_fault_flags[717]          =   1'b0;
assign   tb_i_rf_static_aad_length[717]       =   64'h0000000000000100;
assign   tb_i_aad[717]                        =   tb_i_aad[716];
assign   tb_i_rf_static_plaintext_length[717] =   64'h0000000000000280;
assign   tb_i_plaintext[717]                  =   tb_i_plaintext[716];
assign   tb_o_valid[717]                      =   1'b0;
assign   tb_o_sop[717]                        =   1'b0;
assign   tb_o_ciphertext[717]                 =   tb_o_ciphertext[716];
assign   tb_o_tag_ready[717]                  =   1'b0;
assign   tb_o_tag[717]                        =   tb_o_tag[716];

// CLK no. 718/1240
// *************************************************
assign   tb_i_valid[718]                      =   1'b0;
assign   tb_i_reset[718]                      =   1'b0;
assign   tb_i_sop[718]                        =   1'b0;
assign   tb_i_key_update[718]                 =   1'b0;
assign   tb_i_key[718]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[718]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[718]               =   1'b0;
assign   tb_i_rf_static_encrypt[718]          =   1'b1;
assign   tb_i_clear_fault_flags[718]          =   1'b0;
assign   tb_i_rf_static_aad_length[718]       =   64'h0000000000000100;
assign   tb_i_aad[718]                        =   tb_i_aad[717];
assign   tb_i_rf_static_plaintext_length[718] =   64'h0000000000000280;
assign   tb_i_plaintext[718]                  =   tb_i_plaintext[717];
assign   tb_o_valid[718]                      =   1'b0;
assign   tb_o_sop[718]                        =   1'b0;
assign   tb_o_ciphertext[718]                 =   tb_o_ciphertext[717];
assign   tb_o_tag_ready[718]                  =   1'b0;
assign   tb_o_tag[718]                        =   tb_o_tag[717];

// CLK no. 719/1240
// *************************************************
assign   tb_i_valid[719]                      =   1'b0;
assign   tb_i_reset[719]                      =   1'b0;
assign   tb_i_sop[719]                        =   1'b0;
assign   tb_i_key_update[719]                 =   1'b0;
assign   tb_i_key[719]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[719]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[719]               =   1'b0;
assign   tb_i_rf_static_encrypt[719]          =   1'b1;
assign   tb_i_clear_fault_flags[719]          =   1'b0;
assign   tb_i_rf_static_aad_length[719]       =   64'h0000000000000100;
assign   tb_i_aad[719]                        =   tb_i_aad[718];
assign   tb_i_rf_static_plaintext_length[719] =   64'h0000000000000280;
assign   tb_i_plaintext[719]                  =   tb_i_plaintext[718];
assign   tb_o_valid[719]                      =   1'b0;
assign   tb_o_sop[719]                        =   1'b0;
assign   tb_o_ciphertext[719]                 =   tb_o_ciphertext[718];
assign   tb_o_tag_ready[719]                  =   1'b0;
assign   tb_o_tag[719]                        =   tb_o_tag[718];

// CLK no. 720/1240
// *************************************************
assign   tb_i_valid[720]                      =   1'b0;
assign   tb_i_reset[720]                      =   1'b0;
assign   tb_i_sop[720]                        =   1'b0;
assign   tb_i_key_update[720]                 =   1'b0;
assign   tb_i_key[720]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[720]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[720]               =   1'b0;
assign   tb_i_rf_static_encrypt[720]          =   1'b1;
assign   tb_i_clear_fault_flags[720]          =   1'b0;
assign   tb_i_rf_static_aad_length[720]       =   64'h0000000000000100;
assign   tb_i_aad[720]                        =   tb_i_aad[719];
assign   tb_i_rf_static_plaintext_length[720] =   64'h0000000000000280;
assign   tb_i_plaintext[720]                  =   tb_i_plaintext[719];
assign   tb_o_valid[720]                      =   1'b0;
assign   tb_o_sop[720]                        =   1'b0;
assign   tb_o_ciphertext[720]                 =   tb_o_ciphertext[719];
assign   tb_o_tag_ready[720]                  =   1'b0;
assign   tb_o_tag[720]                        =   tb_o_tag[719];

// CLK no. 721/1240
// *************************************************
assign   tb_i_valid[721]                      =   1'b0;
assign   tb_i_reset[721]                      =   1'b0;
assign   tb_i_sop[721]                        =   1'b0;
assign   tb_i_key_update[721]                 =   1'b0;
assign   tb_i_key[721]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[721]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[721]               =   1'b0;
assign   tb_i_rf_static_encrypt[721]          =   1'b1;
assign   tb_i_clear_fault_flags[721]          =   1'b0;
assign   tb_i_rf_static_aad_length[721]       =   64'h0000000000000100;
assign   tb_i_aad[721]                        =   tb_i_aad[720];
assign   tb_i_rf_static_plaintext_length[721] =   64'h0000000000000280;
assign   tb_i_plaintext[721]                  =   tb_i_plaintext[720];
assign   tb_o_valid[721]                      =   1'b0;
assign   tb_o_sop[721]                        =   1'b0;
assign   tb_o_ciphertext[721]                 =   tb_o_ciphertext[720];
assign   tb_o_tag_ready[721]                  =   1'b0;
assign   tb_o_tag[721]                        =   tb_o_tag[720];

// CLK no. 722/1240
// *************************************************
assign   tb_i_valid[722]                      =   1'b0;
assign   tb_i_reset[722]                      =   1'b0;
assign   tb_i_sop[722]                        =   1'b0;
assign   tb_i_key_update[722]                 =   1'b0;
assign   tb_i_key[722]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[722]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[722]               =   1'b0;
assign   tb_i_rf_static_encrypt[722]          =   1'b1;
assign   tb_i_clear_fault_flags[722]          =   1'b0;
assign   tb_i_rf_static_aad_length[722]       =   64'h0000000000000100;
assign   tb_i_aad[722]                        =   tb_i_aad[721];
assign   tb_i_rf_static_plaintext_length[722] =   64'h0000000000000280;
assign   tb_i_plaintext[722]                  =   tb_i_plaintext[721];
assign   tb_o_valid[722]                      =   1'b0;
assign   tb_o_sop[722]                        =   1'b0;
assign   tb_o_ciphertext[722]                 =   tb_o_ciphertext[721];
assign   tb_o_tag_ready[722]                  =   1'b0;
assign   tb_o_tag[722]                        =   tb_o_tag[721];

// CLK no. 723/1240
// *************************************************
assign   tb_i_valid[723]                      =   1'b0;
assign   tb_i_reset[723]                      =   1'b0;
assign   tb_i_sop[723]                        =   1'b0;
assign   tb_i_key_update[723]                 =   1'b0;
assign   tb_i_key[723]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[723]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[723]               =   1'b0;
assign   tb_i_rf_static_encrypt[723]          =   1'b1;
assign   tb_i_clear_fault_flags[723]          =   1'b0;
assign   tb_i_rf_static_aad_length[723]       =   64'h0000000000000100;
assign   tb_i_aad[723]                        =   tb_i_aad[722];
assign   tb_i_rf_static_plaintext_length[723] =   64'h0000000000000280;
assign   tb_i_plaintext[723]                  =   tb_i_plaintext[722];
assign   tb_o_valid[723]                      =   1'b0;
assign   tb_o_sop[723]                        =   1'b0;
assign   tb_o_ciphertext[723]                 =   tb_o_ciphertext[722];
assign   tb_o_tag_ready[723]                  =   1'b0;
assign   tb_o_tag[723]                        =   tb_o_tag[722];

// CLK no. 724/1240
// *************************************************
assign   tb_i_valid[724]                      =   1'b0;
assign   tb_i_reset[724]                      =   1'b0;
assign   tb_i_sop[724]                        =   1'b0;
assign   tb_i_key_update[724]                 =   1'b0;
assign   tb_i_key[724]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[724]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[724]               =   1'b0;
assign   tb_i_rf_static_encrypt[724]          =   1'b1;
assign   tb_i_clear_fault_flags[724]          =   1'b0;
assign   tb_i_rf_static_aad_length[724]       =   64'h0000000000000100;
assign   tb_i_aad[724]                        =   tb_i_aad[723];
assign   tb_i_rf_static_plaintext_length[724] =   64'h0000000000000280;
assign   tb_i_plaintext[724]                  =   tb_i_plaintext[723];
assign   tb_o_valid[724]                      =   1'b0;
assign   tb_o_sop[724]                        =   1'b0;
assign   tb_o_ciphertext[724]                 =   tb_o_ciphertext[723];
assign   tb_o_tag_ready[724]                  =   1'b0;
assign   tb_o_tag[724]                        =   tb_o_tag[723];

// CLK no. 725/1240
// *************************************************
assign   tb_i_valid[725]                      =   1'b0;
assign   tb_i_reset[725]                      =   1'b0;
assign   tb_i_sop[725]                        =   1'b0;
assign   tb_i_key_update[725]                 =   1'b0;
assign   tb_i_key[725]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[725]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[725]               =   1'b0;
assign   tb_i_rf_static_encrypt[725]          =   1'b1;
assign   tb_i_clear_fault_flags[725]          =   1'b0;
assign   tb_i_rf_static_aad_length[725]       =   64'h0000000000000100;
assign   tb_i_aad[725]                        =   tb_i_aad[724];
assign   tb_i_rf_static_plaintext_length[725] =   64'h0000000000000280;
assign   tb_i_plaintext[725]                  =   tb_i_plaintext[724];
assign   tb_o_valid[725]                      =   1'b0;
assign   tb_o_sop[725]                        =   1'b0;
assign   tb_o_ciphertext[725]                 =   tb_o_ciphertext[724];
assign   tb_o_tag_ready[725]                  =   1'b0;
assign   tb_o_tag[725]                        =   tb_o_tag[724];

// CLK no. 726/1240
// *************************************************
assign   tb_i_valid[726]                      =   1'b0;
assign   tb_i_reset[726]                      =   1'b0;
assign   tb_i_sop[726]                        =   1'b0;
assign   tb_i_key_update[726]                 =   1'b0;
assign   tb_i_key[726]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[726]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[726]               =   1'b0;
assign   tb_i_rf_static_encrypt[726]          =   1'b1;
assign   tb_i_clear_fault_flags[726]          =   1'b0;
assign   tb_i_rf_static_aad_length[726]       =   64'h0000000000000100;
assign   tb_i_aad[726]                        =   tb_i_aad[725];
assign   tb_i_rf_static_plaintext_length[726] =   64'h0000000000000280;
assign   tb_i_plaintext[726]                  =   tb_i_plaintext[725];
assign   tb_o_valid[726]                      =   1'b0;
assign   tb_o_sop[726]                        =   1'b0;
assign   tb_o_ciphertext[726]                 =   tb_o_ciphertext[725];
assign   tb_o_tag_ready[726]                  =   1'b0;
assign   tb_o_tag[726]                        =   tb_o_tag[725];

// CLK no. 727/1240
// *************************************************
assign   tb_i_valid[727]                      =   1'b0;
assign   tb_i_reset[727]                      =   1'b0;
assign   tb_i_sop[727]                        =   1'b0;
assign   tb_i_key_update[727]                 =   1'b0;
assign   tb_i_key[727]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[727]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[727]               =   1'b0;
assign   tb_i_rf_static_encrypt[727]          =   1'b1;
assign   tb_i_clear_fault_flags[727]          =   1'b0;
assign   tb_i_rf_static_aad_length[727]       =   64'h0000000000000100;
assign   tb_i_aad[727]                        =   tb_i_aad[726];
assign   tb_i_rf_static_plaintext_length[727] =   64'h0000000000000280;
assign   tb_i_plaintext[727]                  =   tb_i_plaintext[726];
assign   tb_o_valid[727]                      =   1'b0;
assign   tb_o_sop[727]                        =   1'b0;
assign   tb_o_ciphertext[727]                 =   tb_o_ciphertext[726];
assign   tb_o_tag_ready[727]                  =   1'b0;
assign   tb_o_tag[727]                        =   tb_o_tag[726];

// CLK no. 728/1240
// *************************************************
assign   tb_i_valid[728]                      =   1'b0;
assign   tb_i_reset[728]                      =   1'b0;
assign   tb_i_sop[728]                        =   1'b0;
assign   tb_i_key_update[728]                 =   1'b0;
assign   tb_i_key[728]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[728]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[728]               =   1'b0;
assign   tb_i_rf_static_encrypt[728]          =   1'b1;
assign   tb_i_clear_fault_flags[728]          =   1'b0;
assign   tb_i_rf_static_aad_length[728]       =   64'h0000000000000100;
assign   tb_i_aad[728]                        =   tb_i_aad[727];
assign   tb_i_rf_static_plaintext_length[728] =   64'h0000000000000280;
assign   tb_i_plaintext[728]                  =   tb_i_plaintext[727];
assign   tb_o_valid[728]                      =   1'b0;
assign   tb_o_sop[728]                        =   1'b0;
assign   tb_o_ciphertext[728]                 =   tb_o_ciphertext[727];
assign   tb_o_tag_ready[728]                  =   1'b0;
assign   tb_o_tag[728]                        =   tb_o_tag[727];

// CLK no. 729/1240
// *************************************************
assign   tb_i_valid[729]                      =   1'b0;
assign   tb_i_reset[729]                      =   1'b0;
assign   tb_i_sop[729]                        =   1'b0;
assign   tb_i_key_update[729]                 =   1'b0;
assign   tb_i_key[729]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[729]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[729]               =   1'b0;
assign   tb_i_rf_static_encrypt[729]          =   1'b1;
assign   tb_i_clear_fault_flags[729]          =   1'b0;
assign   tb_i_rf_static_aad_length[729]       =   64'h0000000000000100;
assign   tb_i_aad[729]                        =   tb_i_aad[728];
assign   tb_i_rf_static_plaintext_length[729] =   64'h0000000000000280;
assign   tb_i_plaintext[729]                  =   tb_i_plaintext[728];
assign   tb_o_valid[729]                      =   1'b0;
assign   tb_o_sop[729]                        =   1'b0;
assign   tb_o_ciphertext[729]                 =   tb_o_ciphertext[728];
assign   tb_o_tag_ready[729]                  =   1'b0;
assign   tb_o_tag[729]                        =   tb_o_tag[728];

// CLK no. 730/1240
// *************************************************
assign   tb_i_valid[730]                      =   1'b0;
assign   tb_i_reset[730]                      =   1'b0;
assign   tb_i_sop[730]                        =   1'b0;
assign   tb_i_key_update[730]                 =   1'b0;
assign   tb_i_key[730]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[730]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[730]               =   1'b0;
assign   tb_i_rf_static_encrypt[730]          =   1'b1;
assign   tb_i_clear_fault_flags[730]          =   1'b0;
assign   tb_i_rf_static_aad_length[730]       =   64'h0000000000000100;
assign   tb_i_aad[730]                        =   tb_i_aad[729];
assign   tb_i_rf_static_plaintext_length[730] =   64'h0000000000000280;
assign   tb_i_plaintext[730]                  =   tb_i_plaintext[729];
assign   tb_o_valid[730]                      =   1'b0;
assign   tb_o_sop[730]                        =   1'b0;
assign   tb_o_ciphertext[730]                 =   tb_o_ciphertext[729];
assign   tb_o_tag_ready[730]                  =   1'b0;
assign   tb_o_tag[730]                        =   tb_o_tag[729];

// CLK no. 731/1240
// *************************************************
assign   tb_i_valid[731]                      =   1'b0;
assign   tb_i_reset[731]                      =   1'b0;
assign   tb_i_sop[731]                        =   1'b0;
assign   tb_i_key_update[731]                 =   1'b0;
assign   tb_i_key[731]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[731]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[731]               =   1'b0;
assign   tb_i_rf_static_encrypt[731]          =   1'b1;
assign   tb_i_clear_fault_flags[731]          =   1'b0;
assign   tb_i_rf_static_aad_length[731]       =   64'h0000000000000100;
assign   tb_i_aad[731]                        =   tb_i_aad[730];
assign   tb_i_rf_static_plaintext_length[731] =   64'h0000000000000280;
assign   tb_i_plaintext[731]                  =   tb_i_plaintext[730];
assign   tb_o_valid[731]                      =   1'b0;
assign   tb_o_sop[731]                        =   1'b0;
assign   tb_o_ciphertext[731]                 =   tb_o_ciphertext[730];
assign   tb_o_tag_ready[731]                  =   1'b0;
assign   tb_o_tag[731]                        =   tb_o_tag[730];

// CLK no. 732/1240
// *************************************************
assign   tb_i_valid[732]                      =   1'b0;
assign   tb_i_reset[732]                      =   1'b0;
assign   tb_i_sop[732]                        =   1'b0;
assign   tb_i_key_update[732]                 =   1'b0;
assign   tb_i_key[732]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[732]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[732]               =   1'b0;
assign   tb_i_rf_static_encrypt[732]          =   1'b1;
assign   tb_i_clear_fault_flags[732]          =   1'b0;
assign   tb_i_rf_static_aad_length[732]       =   64'h0000000000000100;
assign   tb_i_aad[732]                        =   tb_i_aad[731];
assign   tb_i_rf_static_plaintext_length[732] =   64'h0000000000000280;
assign   tb_i_plaintext[732]                  =   tb_i_plaintext[731];
assign   tb_o_valid[732]                      =   1'b0;
assign   tb_o_sop[732]                        =   1'b0;
assign   tb_o_ciphertext[732]                 =   tb_o_ciphertext[731];
assign   tb_o_tag_ready[732]                  =   1'b0;
assign   tb_o_tag[732]                        =   tb_o_tag[731];

// CLK no. 733/1240
// *************************************************
assign   tb_i_valid[733]                      =   1'b0;
assign   tb_i_reset[733]                      =   1'b0;
assign   tb_i_sop[733]                        =   1'b0;
assign   tb_i_key_update[733]                 =   1'b0;
assign   tb_i_key[733]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[733]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[733]               =   1'b0;
assign   tb_i_rf_static_encrypt[733]          =   1'b1;
assign   tb_i_clear_fault_flags[733]          =   1'b0;
assign   tb_i_rf_static_aad_length[733]       =   64'h0000000000000100;
assign   tb_i_aad[733]                        =   tb_i_aad[732];
assign   tb_i_rf_static_plaintext_length[733] =   64'h0000000000000280;
assign   tb_i_plaintext[733]                  =   tb_i_plaintext[732];
assign   tb_o_valid[733]                      =   1'b0;
assign   tb_o_sop[733]                        =   1'b0;
assign   tb_o_ciphertext[733]                 =   tb_o_ciphertext[732];
assign   tb_o_tag_ready[733]                  =   1'b0;
assign   tb_o_tag[733]                        =   tb_o_tag[732];

// CLK no. 734/1240
// *************************************************
assign   tb_i_valid[734]                      =   1'b0;
assign   tb_i_reset[734]                      =   1'b0;
assign   tb_i_sop[734]                        =   1'b0;
assign   tb_i_key_update[734]                 =   1'b0;
assign   tb_i_key[734]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[734]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[734]               =   1'b0;
assign   tb_i_rf_static_encrypt[734]          =   1'b1;
assign   tb_i_clear_fault_flags[734]          =   1'b0;
assign   tb_i_rf_static_aad_length[734]       =   64'h0000000000000100;
assign   tb_i_aad[734]                        =   tb_i_aad[733];
assign   tb_i_rf_static_plaintext_length[734] =   64'h0000000000000280;
assign   tb_i_plaintext[734]                  =   tb_i_plaintext[733];
assign   tb_o_valid[734]                      =   1'b0;
assign   tb_o_sop[734]                        =   1'b0;
assign   tb_o_ciphertext[734]                 =   tb_o_ciphertext[733];
assign   tb_o_tag_ready[734]                  =   1'b0;
assign   tb_o_tag[734]                        =   tb_o_tag[733];

// CLK no. 735/1240
// *************************************************
assign   tb_i_valid[735]                      =   1'b0;
assign   tb_i_reset[735]                      =   1'b0;
assign   tb_i_sop[735]                        =   1'b0;
assign   tb_i_key_update[735]                 =   1'b0;
assign   tb_i_key[735]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[735]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[735]               =   1'b0;
assign   tb_i_rf_static_encrypt[735]          =   1'b1;
assign   tb_i_clear_fault_flags[735]          =   1'b0;
assign   tb_i_rf_static_aad_length[735]       =   64'h0000000000000100;
assign   tb_i_aad[735]                        =   tb_i_aad[734];
assign   tb_i_rf_static_plaintext_length[735] =   64'h0000000000000280;
assign   tb_i_plaintext[735]                  =   tb_i_plaintext[734];
assign   tb_o_valid[735]                      =   1'b0;
assign   tb_o_sop[735]                        =   1'b0;
assign   tb_o_ciphertext[735]                 =   tb_o_ciphertext[734];
assign   tb_o_tag_ready[735]                  =   1'b0;
assign   tb_o_tag[735]                        =   tb_o_tag[734];

// CLK no. 736/1240
// *************************************************
assign   tb_i_valid[736]                      =   1'b0;
assign   tb_i_reset[736]                      =   1'b0;
assign   tb_i_sop[736]                        =   1'b0;
assign   tb_i_key_update[736]                 =   1'b0;
assign   tb_i_key[736]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[736]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[736]               =   1'b0;
assign   tb_i_rf_static_encrypt[736]          =   1'b1;
assign   tb_i_clear_fault_flags[736]          =   1'b0;
assign   tb_i_rf_static_aad_length[736]       =   64'h0000000000000100;
assign   tb_i_aad[736]                        =   tb_i_aad[735];
assign   tb_i_rf_static_plaintext_length[736] =   64'h0000000000000280;
assign   tb_i_plaintext[736]                  =   tb_i_plaintext[735];
assign   tb_o_valid[736]                      =   1'b0;
assign   tb_o_sop[736]                        =   1'b0;
assign   tb_o_ciphertext[736]                 =   tb_o_ciphertext[735];
assign   tb_o_tag_ready[736]                  =   1'b0;
assign   tb_o_tag[736]                        =   tb_o_tag[735];

// CLK no. 737/1240
// *************************************************
assign   tb_i_valid[737]                      =   1'b0;
assign   tb_i_reset[737]                      =   1'b0;
assign   tb_i_sop[737]                        =   1'b0;
assign   tb_i_key_update[737]                 =   1'b0;
assign   tb_i_key[737]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[737]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[737]               =   1'b0;
assign   tb_i_rf_static_encrypt[737]          =   1'b1;
assign   tb_i_clear_fault_flags[737]          =   1'b0;
assign   tb_i_rf_static_aad_length[737]       =   64'h0000000000000100;
assign   tb_i_aad[737]                        =   tb_i_aad[736];
assign   tb_i_rf_static_plaintext_length[737] =   64'h0000000000000280;
assign   tb_i_plaintext[737]                  =   tb_i_plaintext[736];
assign   tb_o_valid[737]                      =   1'b0;
assign   tb_o_sop[737]                        =   1'b0;
assign   tb_o_ciphertext[737]                 =   tb_o_ciphertext[736];
assign   tb_o_tag_ready[737]                  =   1'b0;
assign   tb_o_tag[737]                        =   tb_o_tag[736];

// CLK no. 738/1240
// *************************************************
assign   tb_i_valid[738]                      =   1'b0;
assign   tb_i_reset[738]                      =   1'b0;
assign   tb_i_sop[738]                        =   1'b0;
assign   tb_i_key_update[738]                 =   1'b0;
assign   tb_i_key[738]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[738]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[738]               =   1'b0;
assign   tb_i_rf_static_encrypt[738]          =   1'b1;
assign   tb_i_clear_fault_flags[738]          =   1'b0;
assign   tb_i_rf_static_aad_length[738]       =   64'h0000000000000100;
assign   tb_i_aad[738]                        =   tb_i_aad[737];
assign   tb_i_rf_static_plaintext_length[738] =   64'h0000000000000280;
assign   tb_i_plaintext[738]                  =   tb_i_plaintext[737];
assign   tb_o_valid[738]                      =   1'b0;
assign   tb_o_sop[738]                        =   1'b0;
assign   tb_o_ciphertext[738]                 =   tb_o_ciphertext[737];
assign   tb_o_tag_ready[738]                  =   1'b0;
assign   tb_o_tag[738]                        =   tb_o_tag[737];

// CLK no. 739/1240
// *************************************************
assign   tb_i_valid[739]                      =   1'b0;
assign   tb_i_reset[739]                      =   1'b0;
assign   tb_i_sop[739]                        =   1'b0;
assign   tb_i_key_update[739]                 =   1'b0;
assign   tb_i_key[739]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[739]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[739]               =   1'b0;
assign   tb_i_rf_static_encrypt[739]          =   1'b1;
assign   tb_i_clear_fault_flags[739]          =   1'b0;
assign   tb_i_rf_static_aad_length[739]       =   64'h0000000000000100;
assign   tb_i_aad[739]                        =   tb_i_aad[738];
assign   tb_i_rf_static_plaintext_length[739] =   64'h0000000000000280;
assign   tb_i_plaintext[739]                  =   tb_i_plaintext[738];
assign   tb_o_valid[739]                      =   1'b0;
assign   tb_o_sop[739]                        =   1'b0;
assign   tb_o_ciphertext[739]                 =   tb_o_ciphertext[738];
assign   tb_o_tag_ready[739]                  =   1'b0;
assign   tb_o_tag[739]                        =   tb_o_tag[738];

// CLK no. 740/1240
// *************************************************
assign   tb_i_valid[740]                      =   1'b0;
assign   tb_i_reset[740]                      =   1'b0;
assign   tb_i_sop[740]                        =   1'b0;
assign   tb_i_key_update[740]                 =   1'b0;
assign   tb_i_key[740]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[740]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[740]               =   1'b0;
assign   tb_i_rf_static_encrypt[740]          =   1'b1;
assign   tb_i_clear_fault_flags[740]          =   1'b0;
assign   tb_i_rf_static_aad_length[740]       =   64'h0000000000000100;
assign   tb_i_aad[740]                        =   tb_i_aad[739];
assign   tb_i_rf_static_plaintext_length[740] =   64'h0000000000000280;
assign   tb_i_plaintext[740]                  =   tb_i_plaintext[739];
assign   tb_o_valid[740]                      =   1'b0;
assign   tb_o_sop[740]                        =   1'b0;
assign   tb_o_ciphertext[740]                 =   tb_o_ciphertext[739];
assign   tb_o_tag_ready[740]                  =   1'b0;
assign   tb_o_tag[740]                        =   tb_o_tag[739];

// CLK no. 741/1240
// *************************************************
assign   tb_i_valid[741]                      =   1'b0;
assign   tb_i_reset[741]                      =   1'b0;
assign   tb_i_sop[741]                        =   1'b0;
assign   tb_i_key_update[741]                 =   1'b0;
assign   tb_i_key[741]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[741]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[741]               =   1'b0;
assign   tb_i_rf_static_encrypt[741]          =   1'b1;
assign   tb_i_clear_fault_flags[741]          =   1'b0;
assign   tb_i_rf_static_aad_length[741]       =   64'h0000000000000100;
assign   tb_i_aad[741]                        =   tb_i_aad[740];
assign   tb_i_rf_static_plaintext_length[741] =   64'h0000000000000280;
assign   tb_i_plaintext[741]                  =   tb_i_plaintext[740];
assign   tb_o_valid[741]                      =   1'b0;
assign   tb_o_sop[741]                        =   1'b0;
assign   tb_o_ciphertext[741]                 =   tb_o_ciphertext[740];
assign   tb_o_tag_ready[741]                  =   1'b0;
assign   tb_o_tag[741]                        =   tb_o_tag[740];

// CLK no. 742/1240
// *************************************************
assign   tb_i_valid[742]                      =   1'b0;
assign   tb_i_reset[742]                      =   1'b0;
assign   tb_i_sop[742]                        =   1'b0;
assign   tb_i_key_update[742]                 =   1'b0;
assign   tb_i_key[742]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[742]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[742]               =   1'b0;
assign   tb_i_rf_static_encrypt[742]          =   1'b1;
assign   tb_i_clear_fault_flags[742]          =   1'b0;
assign   tb_i_rf_static_aad_length[742]       =   64'h0000000000000100;
assign   tb_i_aad[742]                        =   tb_i_aad[741];
assign   tb_i_rf_static_plaintext_length[742] =   64'h0000000000000280;
assign   tb_i_plaintext[742]                  =   tb_i_plaintext[741];
assign   tb_o_valid[742]                      =   1'b0;
assign   tb_o_sop[742]                        =   1'b0;
assign   tb_o_ciphertext[742]                 =   tb_o_ciphertext[741];
assign   tb_o_tag_ready[742]                  =   1'b0;
assign   tb_o_tag[742]                        =   tb_o_tag[741];

// CLK no. 743/1240
// *************************************************
assign   tb_i_valid[743]                      =   1'b0;
assign   tb_i_reset[743]                      =   1'b0;
assign   tb_i_sop[743]                        =   1'b0;
assign   tb_i_key_update[743]                 =   1'b0;
assign   tb_i_key[743]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[743]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[743]               =   1'b0;
assign   tb_i_rf_static_encrypt[743]          =   1'b1;
assign   tb_i_clear_fault_flags[743]          =   1'b0;
assign   tb_i_rf_static_aad_length[743]       =   64'h0000000000000100;
assign   tb_i_aad[743]                        =   tb_i_aad[742];
assign   tb_i_rf_static_plaintext_length[743] =   64'h0000000000000280;
assign   tb_i_plaintext[743]                  =   tb_i_plaintext[742];
assign   tb_o_valid[743]                      =   1'b0;
assign   tb_o_sop[743]                        =   1'b0;
assign   tb_o_ciphertext[743]                 =   tb_o_ciphertext[742];
assign   tb_o_tag_ready[743]                  =   1'b0;
assign   tb_o_tag[743]                        =   tb_o_tag[742];

// CLK no. 744/1240
// *************************************************
assign   tb_i_valid[744]                      =   1'b0;
assign   tb_i_reset[744]                      =   1'b0;
assign   tb_i_sop[744]                        =   1'b0;
assign   tb_i_key_update[744]                 =   1'b0;
assign   tb_i_key[744]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[744]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[744]               =   1'b0;
assign   tb_i_rf_static_encrypt[744]          =   1'b1;
assign   tb_i_clear_fault_flags[744]          =   1'b0;
assign   tb_i_rf_static_aad_length[744]       =   64'h0000000000000100;
assign   tb_i_aad[744]                        =   tb_i_aad[743];
assign   tb_i_rf_static_plaintext_length[744] =   64'h0000000000000280;
assign   tb_i_plaintext[744]                  =   tb_i_plaintext[743];
assign   tb_o_valid[744]                      =   1'b0;
assign   tb_o_sop[744]                        =   1'b0;
assign   tb_o_ciphertext[744]                 =   tb_o_ciphertext[743];
assign   tb_o_tag_ready[744]                  =   1'b0;
assign   tb_o_tag[744]                        =   tb_o_tag[743];

// CLK no. 745/1240
// *************************************************
assign   tb_i_valid[745]                      =   1'b0;
assign   tb_i_reset[745]                      =   1'b0;
assign   tb_i_sop[745]                        =   1'b0;
assign   tb_i_key_update[745]                 =   1'b0;
assign   tb_i_key[745]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[745]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[745]               =   1'b0;
assign   tb_i_rf_static_encrypt[745]          =   1'b1;
assign   tb_i_clear_fault_flags[745]          =   1'b0;
assign   tb_i_rf_static_aad_length[745]       =   64'h0000000000000100;
assign   tb_i_aad[745]                        =   tb_i_aad[744];
assign   tb_i_rf_static_plaintext_length[745] =   64'h0000000000000280;
assign   tb_i_plaintext[745]                  =   tb_i_plaintext[744];
assign   tb_o_valid[745]                      =   1'b0;
assign   tb_o_sop[745]                        =   1'b0;
assign   tb_o_ciphertext[745]                 =   tb_o_ciphertext[744];
assign   tb_o_tag_ready[745]                  =   1'b0;
assign   tb_o_tag[745]                        =   tb_o_tag[744];

// CLK no. 746/1240
// *************************************************
assign   tb_i_valid[746]                      =   1'b0;
assign   tb_i_reset[746]                      =   1'b0;
assign   tb_i_sop[746]                        =   1'b0;
assign   tb_i_key_update[746]                 =   1'b0;
assign   tb_i_key[746]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[746]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[746]               =   1'b0;
assign   tb_i_rf_static_encrypt[746]          =   1'b1;
assign   tb_i_clear_fault_flags[746]          =   1'b0;
assign   tb_i_rf_static_aad_length[746]       =   64'h0000000000000100;
assign   tb_i_aad[746]                        =   tb_i_aad[745];
assign   tb_i_rf_static_plaintext_length[746] =   64'h0000000000000280;
assign   tb_i_plaintext[746]                  =   tb_i_plaintext[745];
assign   tb_o_valid[746]                      =   1'b0;
assign   tb_o_sop[746]                        =   1'b0;
assign   tb_o_ciphertext[746]                 =   tb_o_ciphertext[745];
assign   tb_o_tag_ready[746]                  =   1'b0;
assign   tb_o_tag[746]                        =   tb_o_tag[745];

// CLK no. 747/1240
// *************************************************
assign   tb_i_valid[747]                      =   1'b0;
assign   tb_i_reset[747]                      =   1'b0;
assign   tb_i_sop[747]                        =   1'b0;
assign   tb_i_key_update[747]                 =   1'b0;
assign   tb_i_key[747]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[747]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[747]               =   1'b0;
assign   tb_i_rf_static_encrypt[747]          =   1'b1;
assign   tb_i_clear_fault_flags[747]          =   1'b0;
assign   tb_i_rf_static_aad_length[747]       =   64'h0000000000000100;
assign   tb_i_aad[747]                        =   tb_i_aad[746];
assign   tb_i_rf_static_plaintext_length[747] =   64'h0000000000000280;
assign   tb_i_plaintext[747]                  =   tb_i_plaintext[746];
assign   tb_o_valid[747]                      =   1'b0;
assign   tb_o_sop[747]                        =   1'b0;
assign   tb_o_ciphertext[747]                 =   tb_o_ciphertext[746];
assign   tb_o_tag_ready[747]                  =   1'b0;
assign   tb_o_tag[747]                        =   tb_o_tag[746];

// CLK no. 748/1240
// *************************************************
assign   tb_i_valid[748]                      =   1'b0;
assign   tb_i_reset[748]                      =   1'b0;
assign   tb_i_sop[748]                        =   1'b0;
assign   tb_i_key_update[748]                 =   1'b0;
assign   tb_i_key[748]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[748]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[748]               =   1'b0;
assign   tb_i_rf_static_encrypt[748]          =   1'b1;
assign   tb_i_clear_fault_flags[748]          =   1'b0;
assign   tb_i_rf_static_aad_length[748]       =   64'h0000000000000100;
assign   tb_i_aad[748]                        =   tb_i_aad[747];
assign   tb_i_rf_static_plaintext_length[748] =   64'h0000000000000280;
assign   tb_i_plaintext[748]                  =   tb_i_plaintext[747];
assign   tb_o_valid[748]                      =   1'b0;
assign   tb_o_sop[748]                        =   1'b0;
assign   tb_o_ciphertext[748]                 =   tb_o_ciphertext[747];
assign   tb_o_tag_ready[748]                  =   1'b0;
assign   tb_o_tag[748]                        =   tb_o_tag[747];

// CLK no. 749/1240
// *************************************************
assign   tb_i_valid[749]                      =   1'b0;
assign   tb_i_reset[749]                      =   1'b0;
assign   tb_i_sop[749]                        =   1'b0;
assign   tb_i_key_update[749]                 =   1'b0;
assign   tb_i_key[749]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[749]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[749]               =   1'b0;
assign   tb_i_rf_static_encrypt[749]          =   1'b1;
assign   tb_i_clear_fault_flags[749]          =   1'b0;
assign   tb_i_rf_static_aad_length[749]       =   64'h0000000000000100;
assign   tb_i_aad[749]                        =   tb_i_aad[748];
assign   tb_i_rf_static_plaintext_length[749] =   64'h0000000000000280;
assign   tb_i_plaintext[749]                  =   tb_i_plaintext[748];
assign   tb_o_valid[749]                      =   1'b0;
assign   tb_o_sop[749]                        =   1'b0;
assign   tb_o_ciphertext[749]                 =   tb_o_ciphertext[748];
assign   tb_o_tag_ready[749]                  =   1'b0;
assign   tb_o_tag[749]                        =   tb_o_tag[748];

// CLK no. 750/1240
// *************************************************
assign   tb_i_valid[750]                      =   1'b0;
assign   tb_i_reset[750]                      =   1'b0;
assign   tb_i_sop[750]                        =   1'b0;
assign   tb_i_key_update[750]                 =   1'b0;
assign   tb_i_key[750]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[750]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[750]               =   1'b0;
assign   tb_i_rf_static_encrypt[750]          =   1'b1;
assign   tb_i_clear_fault_flags[750]          =   1'b0;
assign   tb_i_rf_static_aad_length[750]       =   64'h0000000000000100;
assign   tb_i_aad[750]                        =   tb_i_aad[749];
assign   tb_i_rf_static_plaintext_length[750] =   64'h0000000000000280;
assign   tb_i_plaintext[750]                  =   tb_i_plaintext[749];
assign   tb_o_valid[750]                      =   1'b0;
assign   tb_o_sop[750]                        =   1'b0;
assign   tb_o_ciphertext[750]                 =   tb_o_ciphertext[749];
assign   tb_o_tag_ready[750]                  =   1'b0;
assign   tb_o_tag[750]                        =   tb_o_tag[749];

// CLK no. 751/1240
// *************************************************
assign   tb_i_valid[751]                      =   1'b0;
assign   tb_i_reset[751]                      =   1'b0;
assign   tb_i_sop[751]                        =   1'b0;
assign   tb_i_key_update[751]                 =   1'b0;
assign   tb_i_key[751]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[751]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[751]               =   1'b0;
assign   tb_i_rf_static_encrypt[751]          =   1'b1;
assign   tb_i_clear_fault_flags[751]          =   1'b0;
assign   tb_i_rf_static_aad_length[751]       =   64'h0000000000000100;
assign   tb_i_aad[751]                        =   tb_i_aad[750];
assign   tb_i_rf_static_plaintext_length[751] =   64'h0000000000000280;
assign   tb_i_plaintext[751]                  =   tb_i_plaintext[750];
assign   tb_o_valid[751]                      =   1'b0;
assign   tb_o_sop[751]                        =   1'b0;
assign   tb_o_ciphertext[751]                 =   tb_o_ciphertext[750];
assign   tb_o_tag_ready[751]                  =   1'b0;
assign   tb_o_tag[751]                        =   tb_o_tag[750];

// CLK no. 752/1240
// *************************************************
assign   tb_i_valid[752]                      =   1'b0;
assign   tb_i_reset[752]                      =   1'b0;
assign   tb_i_sop[752]                        =   1'b0;
assign   tb_i_key_update[752]                 =   1'b0;
assign   tb_i_key[752]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[752]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[752]               =   1'b0;
assign   tb_i_rf_static_encrypt[752]          =   1'b1;
assign   tb_i_clear_fault_flags[752]          =   1'b0;
assign   tb_i_rf_static_aad_length[752]       =   64'h0000000000000100;
assign   tb_i_aad[752]                        =   tb_i_aad[751];
assign   tb_i_rf_static_plaintext_length[752] =   64'h0000000000000280;
assign   tb_i_plaintext[752]                  =   tb_i_plaintext[751];
assign   tb_o_valid[752]                      =   1'b0;
assign   tb_o_sop[752]                        =   1'b0;
assign   tb_o_ciphertext[752]                 =   tb_o_ciphertext[751];
assign   tb_o_tag_ready[752]                  =   1'b0;
assign   tb_o_tag[752]                        =   tb_o_tag[751];

// CLK no. 753/1240
// *************************************************
assign   tb_i_valid[753]                      =   1'b0;
assign   tb_i_reset[753]                      =   1'b0;
assign   tb_i_sop[753]                        =   1'b0;
assign   tb_i_key_update[753]                 =   1'b0;
assign   tb_i_key[753]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[753]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[753]               =   1'b0;
assign   tb_i_rf_static_encrypt[753]          =   1'b1;
assign   tb_i_clear_fault_flags[753]          =   1'b0;
assign   tb_i_rf_static_aad_length[753]       =   64'h0000000000000100;
assign   tb_i_aad[753]                        =   tb_i_aad[752];
assign   tb_i_rf_static_plaintext_length[753] =   64'h0000000000000280;
assign   tb_i_plaintext[753]                  =   tb_i_plaintext[752];
assign   tb_o_valid[753]                      =   1'b0;
assign   tb_o_sop[753]                        =   1'b0;
assign   tb_o_ciphertext[753]                 =   tb_o_ciphertext[752];
assign   tb_o_tag_ready[753]                  =   1'b0;
assign   tb_o_tag[753]                        =   tb_o_tag[752];

// CLK no. 754/1240
// *************************************************
assign   tb_i_valid[754]                      =   1'b0;
assign   tb_i_reset[754]                      =   1'b0;
assign   tb_i_sop[754]                        =   1'b0;
assign   tb_i_key_update[754]                 =   1'b0;
assign   tb_i_key[754]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[754]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[754]               =   1'b0;
assign   tb_i_rf_static_encrypt[754]          =   1'b1;
assign   tb_i_clear_fault_flags[754]          =   1'b0;
assign   tb_i_rf_static_aad_length[754]       =   64'h0000000000000100;
assign   tb_i_aad[754]                        =   tb_i_aad[753];
assign   tb_i_rf_static_plaintext_length[754] =   64'h0000000000000280;
assign   tb_i_plaintext[754]                  =   tb_i_plaintext[753];
assign   tb_o_valid[754]                      =   1'b0;
assign   tb_o_sop[754]                        =   1'b0;
assign   tb_o_ciphertext[754]                 =   tb_o_ciphertext[753];
assign   tb_o_tag_ready[754]                  =   1'b0;
assign   tb_o_tag[754]                        =   tb_o_tag[753];

// CLK no. 755/1240
// *************************************************
assign   tb_i_valid[755]                      =   1'b0;
assign   tb_i_reset[755]                      =   1'b0;
assign   tb_i_sop[755]                        =   1'b0;
assign   tb_i_key_update[755]                 =   1'b0;
assign   tb_i_key[755]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[755]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[755]               =   1'b0;
assign   tb_i_rf_static_encrypt[755]          =   1'b1;
assign   tb_i_clear_fault_flags[755]          =   1'b0;
assign   tb_i_rf_static_aad_length[755]       =   64'h0000000000000100;
assign   tb_i_aad[755]                        =   tb_i_aad[754];
assign   tb_i_rf_static_plaintext_length[755] =   64'h0000000000000280;
assign   tb_i_plaintext[755]                  =   tb_i_plaintext[754];
assign   tb_o_valid[755]                      =   1'b1;
assign   tb_o_sop[755]                        =   1'b1;
assign   tb_o_ciphertext[755]                 =   256'h223e5afeebd7c2a7cbb396a3972187090e9422ab31cc11423410c74bacdbd934;
assign   tb_o_tag_ready[755]                  =   1'b0;
assign   tb_o_tag[755]                        =   tb_o_tag[754];

// CLK no. 756/1240
// *************************************************
assign   tb_i_valid[756]                      =   1'b0;
assign   tb_i_reset[756]                      =   1'b0;
assign   tb_i_sop[756]                        =   1'b0;
assign   tb_i_key_update[756]                 =   1'b0;
assign   tb_i_key[756]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[756]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[756]               =   1'b0;
assign   tb_i_rf_static_encrypt[756]          =   1'b1;
assign   tb_i_clear_fault_flags[756]          =   1'b0;
assign   tb_i_rf_static_aad_length[756]       =   64'h0000000000000100;
assign   tb_i_aad[756]                        =   tb_i_aad[755];
assign   tb_i_rf_static_plaintext_length[756] =   64'h0000000000000280;
assign   tb_i_plaintext[756]                  =   tb_i_plaintext[755];
assign   tb_o_valid[756]                      =   1'b1;
assign   tb_o_sop[756]                        =   1'b0;
assign   tb_o_ciphertext[756]                 =   256'h941e51db7769d345ac9b177be96867072fea4d7fb8a6fea6d61dd681c242081d;
assign   tb_o_tag_ready[756]                  =   1'b0;
assign   tb_o_tag[756]                        =   tb_o_tag[755];

// CLK no. 757/1240
// *************************************************
assign   tb_i_valid[757]                      =   1'b0;
assign   tb_i_reset[757]                      =   1'b0;
assign   tb_i_sop[757]                        =   1'b0;
assign   tb_i_key_update[757]                 =   1'b0;
assign   tb_i_key[757]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[757]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[757]               =   1'b0;
assign   tb_i_rf_static_encrypt[757]          =   1'b1;
assign   tb_i_clear_fault_flags[757]          =   1'b0;
assign   tb_i_rf_static_aad_length[757]       =   64'h0000000000000100;
assign   tb_i_aad[757]                        =   tb_i_aad[756];
assign   tb_i_rf_static_plaintext_length[757] =   64'h0000000000000280;
assign   tb_i_plaintext[757]                  =   tb_i_plaintext[756];
assign   tb_o_valid[757]                      =   1'b1;
assign   tb_o_sop[757]                        =   1'b0;
assign   tb_o_ciphertext[757]                 =   256'h4f65dc90187c0a6783f45e910deb1037;
assign   tb_o_tag_ready[757]                  =   1'b0;
assign   tb_o_tag[757]                        =   tb_o_tag[756];

// CLK no. 758/1240
// *************************************************
assign   tb_i_valid[758]                      =   1'b0;
assign   tb_i_reset[758]                      =   1'b0;
assign   tb_i_sop[758]                        =   1'b0;
assign   tb_i_key_update[758]                 =   1'b0;
assign   tb_i_key[758]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[758]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[758]               =   1'b0;
assign   tb_i_rf_static_encrypt[758]          =   1'b1;
assign   tb_i_clear_fault_flags[758]          =   1'b0;
assign   tb_i_rf_static_aad_length[758]       =   64'h0000000000000100;
assign   tb_i_aad[758]                        =   tb_i_aad[757];
assign   tb_i_rf_static_plaintext_length[758] =   64'h0000000000000280;
assign   tb_i_plaintext[758]                  =   tb_i_plaintext[757];
assign   tb_o_valid[758]                      =   1'b0;
assign   tb_o_sop[758]                        =   1'b0;
assign   tb_o_ciphertext[758]                 =   tb_o_ciphertext[757];
assign   tb_o_tag_ready[758]                  =   1'b0;
assign   tb_o_tag[758]                        =   tb_o_tag[757];

// CLK no. 759/1240
// *************************************************
assign   tb_i_valid[759]                      =   1'b0;
assign   tb_i_reset[759]                      =   1'b0;
assign   tb_i_sop[759]                        =   1'b0;
assign   tb_i_key_update[759]                 =   1'b0;
assign   tb_i_key[759]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[759]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[759]               =   1'b0;
assign   tb_i_rf_static_encrypt[759]          =   1'b1;
assign   tb_i_clear_fault_flags[759]          =   1'b0;
assign   tb_i_rf_static_aad_length[759]       =   64'h0000000000000100;
assign   tb_i_aad[759]                        =   tb_i_aad[758];
assign   tb_i_rf_static_plaintext_length[759] =   64'h0000000000000280;
assign   tb_i_plaintext[759]                  =   tb_i_plaintext[758];
assign   tb_o_valid[759]                      =   1'b0;
assign   tb_o_sop[759]                        =   1'b0;
assign   tb_o_ciphertext[759]                 =   tb_o_ciphertext[758];
assign   tb_o_tag_ready[759]                  =   1'b0;
assign   tb_o_tag[759]                        =   tb_o_tag[758];

// CLK no. 760/1240
// *************************************************
assign   tb_i_valid[760]                      =   1'b0;
assign   tb_i_reset[760]                      =   1'b0;
assign   tb_i_sop[760]                        =   1'b0;
assign   tb_i_key_update[760]                 =   1'b0;
assign   tb_i_key[760]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[760]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[760]               =   1'b0;
assign   tb_i_rf_static_encrypt[760]          =   1'b1;
assign   tb_i_clear_fault_flags[760]          =   1'b0;
assign   tb_i_rf_static_aad_length[760]       =   64'h0000000000000100;
assign   tb_i_aad[760]                        =   tb_i_aad[759];
assign   tb_i_rf_static_plaintext_length[760] =   64'h0000000000000280;
assign   tb_i_plaintext[760]                  =   tb_i_plaintext[759];
assign   tb_o_valid[760]                      =   1'b0;
assign   tb_o_sop[760]                        =   1'b0;
assign   tb_o_ciphertext[760]                 =   tb_o_ciphertext[759];
assign   tb_o_tag_ready[760]                  =   1'b0;
assign   tb_o_tag[760]                        =   tb_o_tag[759];

// CLK no. 761/1240
// *************************************************
assign   tb_i_valid[761]                      =   1'b0;
assign   tb_i_reset[761]                      =   1'b0;
assign   tb_i_sop[761]                        =   1'b0;
assign   tb_i_key_update[761]                 =   1'b0;
assign   tb_i_key[761]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[761]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[761]               =   1'b0;
assign   tb_i_rf_static_encrypt[761]          =   1'b1;
assign   tb_i_clear_fault_flags[761]          =   1'b0;
assign   tb_i_rf_static_aad_length[761]       =   64'h0000000000000100;
assign   tb_i_aad[761]                        =   tb_i_aad[760];
assign   tb_i_rf_static_plaintext_length[761] =   64'h0000000000000280;
assign   tb_i_plaintext[761]                  =   tb_i_plaintext[760];
assign   tb_o_valid[761]                      =   1'b0;
assign   tb_o_sop[761]                        =   1'b0;
assign   tb_o_ciphertext[761]                 =   tb_o_ciphertext[760];
assign   tb_o_tag_ready[761]                  =   1'b0;
assign   tb_o_tag[761]                        =   tb_o_tag[760];

// CLK no. 762/1240
// *************************************************
assign   tb_i_valid[762]                      =   1'b0;
assign   tb_i_reset[762]                      =   1'b0;
assign   tb_i_sop[762]                        =   1'b0;
assign   tb_i_key_update[762]                 =   1'b0;
assign   tb_i_key[762]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[762]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[762]               =   1'b0;
assign   tb_i_rf_static_encrypt[762]          =   1'b1;
assign   tb_i_clear_fault_flags[762]          =   1'b0;
assign   tb_i_rf_static_aad_length[762]       =   64'h0000000000000100;
assign   tb_i_aad[762]                        =   tb_i_aad[761];
assign   tb_i_rf_static_plaintext_length[762] =   64'h0000000000000280;
assign   tb_i_plaintext[762]                  =   tb_i_plaintext[761];
assign   tb_o_valid[762]                      =   1'b0;
assign   tb_o_sop[762]                        =   1'b0;
assign   tb_o_ciphertext[762]                 =   tb_o_ciphertext[761];
assign   tb_o_tag_ready[762]                  =   1'b0;
assign   tb_o_tag[762]                        =   tb_o_tag[761];

// CLK no. 763/1240
// *************************************************
assign   tb_i_valid[763]                      =   1'b0;
assign   tb_i_reset[763]                      =   1'b0;
assign   tb_i_sop[763]                        =   1'b0;
assign   tb_i_key_update[763]                 =   1'b0;
assign   tb_i_key[763]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[763]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[763]               =   1'b0;
assign   tb_i_rf_static_encrypt[763]          =   1'b1;
assign   tb_i_clear_fault_flags[763]          =   1'b0;
assign   tb_i_rf_static_aad_length[763]       =   64'h0000000000000100;
assign   tb_i_aad[763]                        =   tb_i_aad[762];
assign   tb_i_rf_static_plaintext_length[763] =   64'h0000000000000280;
assign   tb_i_plaintext[763]                  =   tb_i_plaintext[762];
assign   tb_o_valid[763]                      =   1'b0;
assign   tb_o_sop[763]                        =   1'b0;
assign   tb_o_ciphertext[763]                 =   tb_o_ciphertext[762];
assign   tb_o_tag_ready[763]                  =   1'b0;
assign   tb_o_tag[763]                        =   tb_o_tag[762];

// CLK no. 764/1240
// *************************************************
assign   tb_i_valid[764]                      =   1'b0;
assign   tb_i_reset[764]                      =   1'b0;
assign   tb_i_sop[764]                        =   1'b0;
assign   tb_i_key_update[764]                 =   1'b0;
assign   tb_i_key[764]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[764]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[764]               =   1'b0;
assign   tb_i_rf_static_encrypt[764]          =   1'b1;
assign   tb_i_clear_fault_flags[764]          =   1'b0;
assign   tb_i_rf_static_aad_length[764]       =   64'h0000000000000100;
assign   tb_i_aad[764]                        =   tb_i_aad[763];
assign   tb_i_rf_static_plaintext_length[764] =   64'h0000000000000280;
assign   tb_i_plaintext[764]                  =   tb_i_plaintext[763];
assign   tb_o_valid[764]                      =   1'b0;
assign   tb_o_sop[764]                        =   1'b0;
assign   tb_o_ciphertext[764]                 =   tb_o_ciphertext[763];
assign   tb_o_tag_ready[764]                  =   1'b0;
assign   tb_o_tag[764]                        =   tb_o_tag[763];

// CLK no. 765/1240
// *************************************************
assign   tb_i_valid[765]                      =   1'b0;
assign   tb_i_reset[765]                      =   1'b0;
assign   tb_i_sop[765]                        =   1'b0;
assign   tb_i_key_update[765]                 =   1'b0;
assign   tb_i_key[765]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[765]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[765]               =   1'b0;
assign   tb_i_rf_static_encrypt[765]          =   1'b1;
assign   tb_i_clear_fault_flags[765]          =   1'b0;
assign   tb_i_rf_static_aad_length[765]       =   64'h0000000000000100;
assign   tb_i_aad[765]                        =   tb_i_aad[764];
assign   tb_i_rf_static_plaintext_length[765] =   64'h0000000000000280;
assign   tb_i_plaintext[765]                  =   tb_i_plaintext[764];
assign   tb_o_valid[765]                      =   1'b0;
assign   tb_o_sop[765]                        =   1'b0;
assign   tb_o_ciphertext[765]                 =   tb_o_ciphertext[764];
assign   tb_o_tag_ready[765]                  =   1'b1;
assign   tb_o_tag[765]                        =   128'h59e24d562cb29281010fa6efbd020a48;

// CLK no. 766/1240
// *************************************************
assign   tb_i_valid[766]                      =   1'b0;
assign   tb_i_reset[766]                      =   1'b0;
assign   tb_i_sop[766]                        =   1'b0;
assign   tb_i_key_update[766]                 =   1'b0;
assign   tb_i_key[766]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[766]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[766]               =   1'b0;
assign   tb_i_rf_static_encrypt[766]          =   1'b1;
assign   tb_i_clear_fault_flags[766]          =   1'b0;
assign   tb_i_rf_static_aad_length[766]       =   64'h0000000000000100;
assign   tb_i_aad[766]                        =   tb_i_aad[765];
assign   tb_i_rf_static_plaintext_length[766] =   64'h0000000000000280;
assign   tb_i_plaintext[766]                  =   tb_i_plaintext[765];
assign   tb_o_valid[766]                      =   1'b0;
assign   tb_o_sop[766]                        =   1'b0;
assign   tb_o_ciphertext[766]                 =   tb_o_ciphertext[765];
assign   tb_o_tag_ready[766]                  =   1'b0;
assign   tb_o_tag[766]                        =   tb_o_tag[765];

// CLK no. 767/1240
// *************************************************
assign   tb_i_valid[767]                      =   1'b0;
assign   tb_i_reset[767]                      =   1'b0;
assign   tb_i_sop[767]                        =   1'b0;
assign   tb_i_key_update[767]                 =   1'b0;
assign   tb_i_key[767]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[767]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[767]               =   1'b0;
assign   tb_i_rf_static_encrypt[767]          =   1'b1;
assign   tb_i_clear_fault_flags[767]          =   1'b0;
assign   tb_i_rf_static_aad_length[767]       =   64'h0000000000000100;
assign   tb_i_aad[767]                        =   tb_i_aad[766];
assign   tb_i_rf_static_plaintext_length[767] =   64'h0000000000000280;
assign   tb_i_plaintext[767]                  =   tb_i_plaintext[766];
assign   tb_o_valid[767]                      =   1'b0;
assign   tb_o_sop[767]                        =   1'b0;
assign   tb_o_ciphertext[767]                 =   tb_o_ciphertext[766];
assign   tb_o_tag_ready[767]                  =   1'b0;
assign   tb_o_tag[767]                        =   tb_o_tag[766];

// CLK no. 768/1240
// *************************************************
assign   tb_i_valid[768]                      =   1'b0;
assign   tb_i_reset[768]                      =   1'b0;
assign   tb_i_sop[768]                        =   1'b1;
assign   tb_i_key_update[768]                 =   1'b0;
assign   tb_i_key[768]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[768]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[768]               =   1'b0;
assign   tb_i_rf_static_encrypt[768]          =   1'b1;
assign   tb_i_clear_fault_flags[768]          =   1'b0;
assign   tb_i_rf_static_aad_length[768]       =   64'h0000000000000100;
assign   tb_i_aad[768]                        =   tb_i_aad[767];
assign   tb_i_rf_static_plaintext_length[768] =   64'h0000000000000280;
assign   tb_i_plaintext[768]                  =   tb_i_plaintext[767];
assign   tb_o_valid[768]                      =   1'b0;
assign   tb_o_sop[768]                        =   1'b0;
assign   tb_o_ciphertext[768]                 =   tb_o_ciphertext[767];
assign   tb_o_tag_ready[768]                  =   1'b0;
assign   tb_o_tag[768]                        =   tb_o_tag[767];

// CLK no. 769/1240
// *************************************************
assign   tb_i_valid[769]                      =   1'b1;
assign   tb_i_reset[769]                      =   1'b0;
assign   tb_i_sop[769]                        =   1'b0;
assign   tb_i_key_update[769]                 =   1'b0;
assign   tb_i_key[769]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[769]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[769]               =   1'b0;
assign   tb_i_rf_static_encrypt[769]          =   1'b1;
assign   tb_i_clear_fault_flags[769]          =   1'b0;
assign   tb_i_rf_static_aad_length[769]       =   64'h0000000000000100;
assign   tb_i_aad[769]                        =   256'hb2d726857590280591728d44a4ae8579850cd6135964c678b3a812db6a2296cc;
assign   tb_i_rf_static_plaintext_length[769] =   64'h0000000000000280;
assign   tb_i_plaintext[769]                  =   tb_i_plaintext[768];
assign   tb_o_valid[769]                      =   1'b0;
assign   tb_o_sop[769]                        =   1'b0;
assign   tb_o_ciphertext[769]                 =   tb_o_ciphertext[768];
assign   tb_o_tag_ready[769]                  =   1'b0;
assign   tb_o_tag[769]                        =   tb_o_tag[768];

// CLK no. 770/1240
// *************************************************
assign   tb_i_valid[770]                      =   1'b1;
assign   tb_i_reset[770]                      =   1'b0;
assign   tb_i_sop[770]                        =   1'b0;
assign   tb_i_key_update[770]                 =   1'b0;
assign   tb_i_key[770]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[770]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[770]               =   1'b0;
assign   tb_i_rf_static_encrypt[770]          =   1'b1;
assign   tb_i_clear_fault_flags[770]          =   1'b0;
assign   tb_i_rf_static_aad_length[770]       =   64'h0000000000000100;
assign   tb_i_aad[770]                        =   tb_i_aad[769];
assign   tb_i_rf_static_plaintext_length[770] =   64'h0000000000000280;
assign   tb_i_plaintext[770]                  =   256'hfeaf9e695f6cb2c5bc51c92a36c484e745e92b4ce2309ecbf9279fcdc7b08d47;
assign   tb_o_valid[770]                      =   1'b0;
assign   tb_o_sop[770]                        =   1'b0;
assign   tb_o_ciphertext[770]                 =   tb_o_ciphertext[769];
assign   tb_o_tag_ready[770]                  =   1'b0;
assign   tb_o_tag[770]                        =   tb_o_tag[769];

// CLK no. 771/1240
// *************************************************
assign   tb_i_valid[771]                      =   1'b1;
assign   tb_i_reset[771]                      =   1'b0;
assign   tb_i_sop[771]                        =   1'b0;
assign   tb_i_key_update[771]                 =   1'b0;
assign   tb_i_key[771]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[771]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[771]               =   1'b0;
assign   tb_i_rf_static_encrypt[771]          =   1'b1;
assign   tb_i_clear_fault_flags[771]          =   1'b0;
assign   tb_i_rf_static_aad_length[771]       =   64'h0000000000000100;
assign   tb_i_aad[771]                        =   tb_i_aad[770];
assign   tb_i_rf_static_plaintext_length[771] =   64'h0000000000000280;
assign   tb_i_plaintext[771]                  =   256'h43139f0e6f40ba8f0ab0ce9a5d0c3703db1b6047502a6b094350597e75d3e952;
assign   tb_o_valid[771]                      =   1'b0;
assign   tb_o_sop[771]                        =   1'b0;
assign   tb_o_ciphertext[771]                 =   tb_o_ciphertext[770];
assign   tb_o_tag_ready[771]                  =   1'b0;
assign   tb_o_tag[771]                        =   tb_o_tag[770];

// CLK no. 772/1240
// *************************************************
assign   tb_i_valid[772]                      =   1'b1;
assign   tb_i_reset[772]                      =   1'b0;
assign   tb_i_sop[772]                        =   1'b0;
assign   tb_i_key_update[772]                 =   1'b0;
assign   tb_i_key[772]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[772]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[772]               =   1'b0;
assign   tb_i_rf_static_encrypt[772]          =   1'b1;
assign   tb_i_clear_fault_flags[772]          =   1'b0;
assign   tb_i_rf_static_aad_length[772]       =   64'h0000000000000100;
assign   tb_i_aad[772]                        =   tb_i_aad[771];
assign   tb_i_rf_static_plaintext_length[772] =   64'h0000000000000280;
assign   tb_i_plaintext[772]                  =   256'he06d3d286e1ab8bbd7fa3814a21c2df2;
assign   tb_o_valid[772]                      =   1'b0;
assign   tb_o_sop[772]                        =   1'b0;
assign   tb_o_ciphertext[772]                 =   tb_o_ciphertext[771];
assign   tb_o_tag_ready[772]                  =   1'b0;
assign   tb_o_tag[772]                        =   tb_o_tag[771];

// CLK no. 773/1240
// *************************************************
assign   tb_i_valid[773]                      =   1'b0;
assign   tb_i_reset[773]                      =   1'b0;
assign   tb_i_sop[773]                        =   1'b0;
assign   tb_i_key_update[773]                 =   1'b0;
assign   tb_i_key[773]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[773]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[773]               =   1'b0;
assign   tb_i_rf_static_encrypt[773]          =   1'b1;
assign   tb_i_clear_fault_flags[773]          =   1'b0;
assign   tb_i_rf_static_aad_length[773]       =   64'h0000000000000100;
assign   tb_i_aad[773]                        =   tb_i_aad[772];
assign   tb_i_rf_static_plaintext_length[773] =   64'h0000000000000280;
assign   tb_i_plaintext[773]                  =   tb_i_plaintext[772];
assign   tb_o_valid[773]                      =   1'b0;
assign   tb_o_sop[773]                        =   1'b0;
assign   tb_o_ciphertext[773]                 =   tb_o_ciphertext[772];
assign   tb_o_tag_ready[773]                  =   1'b0;
assign   tb_o_tag[773]                        =   tb_o_tag[772];

// CLK no. 774/1240
// *************************************************
assign   tb_i_valid[774]                      =   1'b0;
assign   tb_i_reset[774]                      =   1'b0;
assign   tb_i_sop[774]                        =   1'b0;
assign   tb_i_key_update[774]                 =   1'b0;
assign   tb_i_key[774]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[774]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[774]               =   1'b0;
assign   tb_i_rf_static_encrypt[774]          =   1'b1;
assign   tb_i_clear_fault_flags[774]          =   1'b0;
assign   tb_i_rf_static_aad_length[774]       =   64'h0000000000000100;
assign   tb_i_aad[774]                        =   tb_i_aad[773];
assign   tb_i_rf_static_plaintext_length[774] =   64'h0000000000000280;
assign   tb_i_plaintext[774]                  =   tb_i_plaintext[773];
assign   tb_o_valid[774]                      =   1'b0;
assign   tb_o_sop[774]                        =   1'b0;
assign   tb_o_ciphertext[774]                 =   tb_o_ciphertext[773];
assign   tb_o_tag_ready[774]                  =   1'b0;
assign   tb_o_tag[774]                        =   tb_o_tag[773];

// CLK no. 775/1240
// *************************************************
assign   tb_i_valid[775]                      =   1'b0;
assign   tb_i_reset[775]                      =   1'b0;
assign   tb_i_sop[775]                        =   1'b0;
assign   tb_i_key_update[775]                 =   1'b0;
assign   tb_i_key[775]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[775]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[775]               =   1'b0;
assign   tb_i_rf_static_encrypt[775]          =   1'b1;
assign   tb_i_clear_fault_flags[775]          =   1'b0;
assign   tb_i_rf_static_aad_length[775]       =   64'h0000000000000100;
assign   tb_i_aad[775]                        =   tb_i_aad[774];
assign   tb_i_rf_static_plaintext_length[775] =   64'h0000000000000280;
assign   tb_i_plaintext[775]                  =   tb_i_plaintext[774];
assign   tb_o_valid[775]                      =   1'b0;
assign   tb_o_sop[775]                        =   1'b0;
assign   tb_o_ciphertext[775]                 =   tb_o_ciphertext[774];
assign   tb_o_tag_ready[775]                  =   1'b0;
assign   tb_o_tag[775]                        =   tb_o_tag[774];

// CLK no. 776/1240
// *************************************************
assign   tb_i_valid[776]                      =   1'b0;
assign   tb_i_reset[776]                      =   1'b0;
assign   tb_i_sop[776]                        =   1'b0;
assign   tb_i_key_update[776]                 =   1'b0;
assign   tb_i_key[776]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[776]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[776]               =   1'b0;
assign   tb_i_rf_static_encrypt[776]          =   1'b1;
assign   tb_i_clear_fault_flags[776]          =   1'b0;
assign   tb_i_rf_static_aad_length[776]       =   64'h0000000000000100;
assign   tb_i_aad[776]                        =   tb_i_aad[775];
assign   tb_i_rf_static_plaintext_length[776] =   64'h0000000000000280;
assign   tb_i_plaintext[776]                  =   tb_i_plaintext[775];
assign   tb_o_valid[776]                      =   1'b0;
assign   tb_o_sop[776]                        =   1'b0;
assign   tb_o_ciphertext[776]                 =   tb_o_ciphertext[775];
assign   tb_o_tag_ready[776]                  =   1'b0;
assign   tb_o_tag[776]                        =   tb_o_tag[775];

// CLK no. 777/1240
// *************************************************
assign   tb_i_valid[777]                      =   1'b0;
assign   tb_i_reset[777]                      =   1'b0;
assign   tb_i_sop[777]                        =   1'b0;
assign   tb_i_key_update[777]                 =   1'b0;
assign   tb_i_key[777]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[777]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[777]               =   1'b0;
assign   tb_i_rf_static_encrypt[777]          =   1'b1;
assign   tb_i_clear_fault_flags[777]          =   1'b0;
assign   tb_i_rf_static_aad_length[777]       =   64'h0000000000000100;
assign   tb_i_aad[777]                        =   tb_i_aad[776];
assign   tb_i_rf_static_plaintext_length[777] =   64'h0000000000000280;
assign   tb_i_plaintext[777]                  =   tb_i_plaintext[776];
assign   tb_o_valid[777]                      =   1'b0;
assign   tb_o_sop[777]                        =   1'b0;
assign   tb_o_ciphertext[777]                 =   tb_o_ciphertext[776];
assign   tb_o_tag_ready[777]                  =   1'b0;
assign   tb_o_tag[777]                        =   tb_o_tag[776];

// CLK no. 778/1240
// *************************************************
assign   tb_i_valid[778]                      =   1'b0;
assign   tb_i_reset[778]                      =   1'b0;
assign   tb_i_sop[778]                        =   1'b0;
assign   tb_i_key_update[778]                 =   1'b0;
assign   tb_i_key[778]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[778]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[778]               =   1'b0;
assign   tb_i_rf_static_encrypt[778]          =   1'b1;
assign   tb_i_clear_fault_flags[778]          =   1'b0;
assign   tb_i_rf_static_aad_length[778]       =   64'h0000000000000100;
assign   tb_i_aad[778]                        =   tb_i_aad[777];
assign   tb_i_rf_static_plaintext_length[778] =   64'h0000000000000280;
assign   tb_i_plaintext[778]                  =   tb_i_plaintext[777];
assign   tb_o_valid[778]                      =   1'b0;
assign   tb_o_sop[778]                        =   1'b0;
assign   tb_o_ciphertext[778]                 =   tb_o_ciphertext[777];
assign   tb_o_tag_ready[778]                  =   1'b0;
assign   tb_o_tag[778]                        =   tb_o_tag[777];

// CLK no. 779/1240
// *************************************************
assign   tb_i_valid[779]                      =   1'b0;
assign   tb_i_reset[779]                      =   1'b0;
assign   tb_i_sop[779]                        =   1'b0;
assign   tb_i_key_update[779]                 =   1'b0;
assign   tb_i_key[779]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[779]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[779]               =   1'b0;
assign   tb_i_rf_static_encrypt[779]          =   1'b1;
assign   tb_i_clear_fault_flags[779]          =   1'b0;
assign   tb_i_rf_static_aad_length[779]       =   64'h0000000000000100;
assign   tb_i_aad[779]                        =   tb_i_aad[778];
assign   tb_i_rf_static_plaintext_length[779] =   64'h0000000000000280;
assign   tb_i_plaintext[779]                  =   tb_i_plaintext[778];
assign   tb_o_valid[779]                      =   1'b0;
assign   tb_o_sop[779]                        =   1'b0;
assign   tb_o_ciphertext[779]                 =   tb_o_ciphertext[778];
assign   tb_o_tag_ready[779]                  =   1'b0;
assign   tb_o_tag[779]                        =   tb_o_tag[778];

// CLK no. 780/1240
// *************************************************
assign   tb_i_valid[780]                      =   1'b0;
assign   tb_i_reset[780]                      =   1'b0;
assign   tb_i_sop[780]                        =   1'b0;
assign   tb_i_key_update[780]                 =   1'b0;
assign   tb_i_key[780]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[780]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[780]               =   1'b0;
assign   tb_i_rf_static_encrypt[780]          =   1'b1;
assign   tb_i_clear_fault_flags[780]          =   1'b0;
assign   tb_i_rf_static_aad_length[780]       =   64'h0000000000000100;
assign   tb_i_aad[780]                        =   tb_i_aad[779];
assign   tb_i_rf_static_plaintext_length[780] =   64'h0000000000000280;
assign   tb_i_plaintext[780]                  =   tb_i_plaintext[779];
assign   tb_o_valid[780]                      =   1'b0;
assign   tb_o_sop[780]                        =   1'b0;
assign   tb_o_ciphertext[780]                 =   tb_o_ciphertext[779];
assign   tb_o_tag_ready[780]                  =   1'b0;
assign   tb_o_tag[780]                        =   tb_o_tag[779];

// CLK no. 781/1240
// *************************************************
assign   tb_i_valid[781]                      =   1'b0;
assign   tb_i_reset[781]                      =   1'b0;
assign   tb_i_sop[781]                        =   1'b0;
assign   tb_i_key_update[781]                 =   1'b0;
assign   tb_i_key[781]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[781]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[781]               =   1'b0;
assign   tb_i_rf_static_encrypt[781]          =   1'b1;
assign   tb_i_clear_fault_flags[781]          =   1'b0;
assign   tb_i_rf_static_aad_length[781]       =   64'h0000000000000100;
assign   tb_i_aad[781]                        =   tb_i_aad[780];
assign   tb_i_rf_static_plaintext_length[781] =   64'h0000000000000280;
assign   tb_i_plaintext[781]                  =   tb_i_plaintext[780];
assign   tb_o_valid[781]                      =   1'b0;
assign   tb_o_sop[781]                        =   1'b0;
assign   tb_o_ciphertext[781]                 =   tb_o_ciphertext[780];
assign   tb_o_tag_ready[781]                  =   1'b0;
assign   tb_o_tag[781]                        =   tb_o_tag[780];

// CLK no. 782/1240
// *************************************************
assign   tb_i_valid[782]                      =   1'b0;
assign   tb_i_reset[782]                      =   1'b0;
assign   tb_i_sop[782]                        =   1'b0;
assign   tb_i_key_update[782]                 =   1'b0;
assign   tb_i_key[782]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[782]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[782]               =   1'b0;
assign   tb_i_rf_static_encrypt[782]          =   1'b1;
assign   tb_i_clear_fault_flags[782]          =   1'b0;
assign   tb_i_rf_static_aad_length[782]       =   64'h0000000000000100;
assign   tb_i_aad[782]                        =   tb_i_aad[781];
assign   tb_i_rf_static_plaintext_length[782] =   64'h0000000000000280;
assign   tb_i_plaintext[782]                  =   tb_i_plaintext[781];
assign   tb_o_valid[782]                      =   1'b0;
assign   tb_o_sop[782]                        =   1'b0;
assign   tb_o_ciphertext[782]                 =   tb_o_ciphertext[781];
assign   tb_o_tag_ready[782]                  =   1'b0;
assign   tb_o_tag[782]                        =   tb_o_tag[781];

// CLK no. 783/1240
// *************************************************
assign   tb_i_valid[783]                      =   1'b0;
assign   tb_i_reset[783]                      =   1'b0;
assign   tb_i_sop[783]                        =   1'b0;
assign   tb_i_key_update[783]                 =   1'b0;
assign   tb_i_key[783]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[783]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[783]               =   1'b0;
assign   tb_i_rf_static_encrypt[783]          =   1'b1;
assign   tb_i_clear_fault_flags[783]          =   1'b0;
assign   tb_i_rf_static_aad_length[783]       =   64'h0000000000000100;
assign   tb_i_aad[783]                        =   tb_i_aad[782];
assign   tb_i_rf_static_plaintext_length[783] =   64'h0000000000000280;
assign   tb_i_plaintext[783]                  =   tb_i_plaintext[782];
assign   tb_o_valid[783]                      =   1'b0;
assign   tb_o_sop[783]                        =   1'b0;
assign   tb_o_ciphertext[783]                 =   tb_o_ciphertext[782];
assign   tb_o_tag_ready[783]                  =   1'b0;
assign   tb_o_tag[783]                        =   tb_o_tag[782];

// CLK no. 784/1240
// *************************************************
assign   tb_i_valid[784]                      =   1'b0;
assign   tb_i_reset[784]                      =   1'b0;
assign   tb_i_sop[784]                        =   1'b0;
assign   tb_i_key_update[784]                 =   1'b0;
assign   tb_i_key[784]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[784]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[784]               =   1'b0;
assign   tb_i_rf_static_encrypt[784]          =   1'b1;
assign   tb_i_clear_fault_flags[784]          =   1'b0;
assign   tb_i_rf_static_aad_length[784]       =   64'h0000000000000100;
assign   tb_i_aad[784]                        =   tb_i_aad[783];
assign   tb_i_rf_static_plaintext_length[784] =   64'h0000000000000280;
assign   tb_i_plaintext[784]                  =   tb_i_plaintext[783];
assign   tb_o_valid[784]                      =   1'b0;
assign   tb_o_sop[784]                        =   1'b0;
assign   tb_o_ciphertext[784]                 =   tb_o_ciphertext[783];
assign   tb_o_tag_ready[784]                  =   1'b0;
assign   tb_o_tag[784]                        =   tb_o_tag[783];

// CLK no. 785/1240
// *************************************************
assign   tb_i_valid[785]                      =   1'b0;
assign   tb_i_reset[785]                      =   1'b0;
assign   tb_i_sop[785]                        =   1'b0;
assign   tb_i_key_update[785]                 =   1'b0;
assign   tb_i_key[785]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[785]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[785]               =   1'b0;
assign   tb_i_rf_static_encrypt[785]          =   1'b1;
assign   tb_i_clear_fault_flags[785]          =   1'b0;
assign   tb_i_rf_static_aad_length[785]       =   64'h0000000000000100;
assign   tb_i_aad[785]                        =   tb_i_aad[784];
assign   tb_i_rf_static_plaintext_length[785] =   64'h0000000000000280;
assign   tb_i_plaintext[785]                  =   tb_i_plaintext[784];
assign   tb_o_valid[785]                      =   1'b0;
assign   tb_o_sop[785]                        =   1'b0;
assign   tb_o_ciphertext[785]                 =   tb_o_ciphertext[784];
assign   tb_o_tag_ready[785]                  =   1'b0;
assign   tb_o_tag[785]                        =   tb_o_tag[784];

// CLK no. 786/1240
// *************************************************
assign   tb_i_valid[786]                      =   1'b0;
assign   tb_i_reset[786]                      =   1'b0;
assign   tb_i_sop[786]                        =   1'b0;
assign   tb_i_key_update[786]                 =   1'b0;
assign   tb_i_key[786]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[786]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[786]               =   1'b0;
assign   tb_i_rf_static_encrypt[786]          =   1'b1;
assign   tb_i_clear_fault_flags[786]          =   1'b0;
assign   tb_i_rf_static_aad_length[786]       =   64'h0000000000000100;
assign   tb_i_aad[786]                        =   tb_i_aad[785];
assign   tb_i_rf_static_plaintext_length[786] =   64'h0000000000000280;
assign   tb_i_plaintext[786]                  =   tb_i_plaintext[785];
assign   tb_o_valid[786]                      =   1'b0;
assign   tb_o_sop[786]                        =   1'b0;
assign   tb_o_ciphertext[786]                 =   tb_o_ciphertext[785];
assign   tb_o_tag_ready[786]                  =   1'b0;
assign   tb_o_tag[786]                        =   tb_o_tag[785];

// CLK no. 787/1240
// *************************************************
assign   tb_i_valid[787]                      =   1'b0;
assign   tb_i_reset[787]                      =   1'b0;
assign   tb_i_sop[787]                        =   1'b0;
assign   tb_i_key_update[787]                 =   1'b0;
assign   tb_i_key[787]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[787]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[787]               =   1'b0;
assign   tb_i_rf_static_encrypt[787]          =   1'b1;
assign   tb_i_clear_fault_flags[787]          =   1'b0;
assign   tb_i_rf_static_aad_length[787]       =   64'h0000000000000100;
assign   tb_i_aad[787]                        =   tb_i_aad[786];
assign   tb_i_rf_static_plaintext_length[787] =   64'h0000000000000280;
assign   tb_i_plaintext[787]                  =   tb_i_plaintext[786];
assign   tb_o_valid[787]                      =   1'b0;
assign   tb_o_sop[787]                        =   1'b0;
assign   tb_o_ciphertext[787]                 =   tb_o_ciphertext[786];
assign   tb_o_tag_ready[787]                  =   1'b0;
assign   tb_o_tag[787]                        =   tb_o_tag[786];

// CLK no. 788/1240
// *************************************************
assign   tb_i_valid[788]                      =   1'b0;
assign   tb_i_reset[788]                      =   1'b0;
assign   tb_i_sop[788]                        =   1'b0;
assign   tb_i_key_update[788]                 =   1'b0;
assign   tb_i_key[788]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[788]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[788]               =   1'b0;
assign   tb_i_rf_static_encrypt[788]          =   1'b1;
assign   tb_i_clear_fault_flags[788]          =   1'b0;
assign   tb_i_rf_static_aad_length[788]       =   64'h0000000000000100;
assign   tb_i_aad[788]                        =   tb_i_aad[787];
assign   tb_i_rf_static_plaintext_length[788] =   64'h0000000000000280;
assign   tb_i_plaintext[788]                  =   tb_i_plaintext[787];
assign   tb_o_valid[788]                      =   1'b0;
assign   tb_o_sop[788]                        =   1'b0;
assign   tb_o_ciphertext[788]                 =   tb_o_ciphertext[787];
assign   tb_o_tag_ready[788]                  =   1'b0;
assign   tb_o_tag[788]                        =   tb_o_tag[787];

// CLK no. 789/1240
// *************************************************
assign   tb_i_valid[789]                      =   1'b0;
assign   tb_i_reset[789]                      =   1'b0;
assign   tb_i_sop[789]                        =   1'b0;
assign   tb_i_key_update[789]                 =   1'b0;
assign   tb_i_key[789]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[789]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[789]               =   1'b0;
assign   tb_i_rf_static_encrypt[789]          =   1'b1;
assign   tb_i_clear_fault_flags[789]          =   1'b0;
assign   tb_i_rf_static_aad_length[789]       =   64'h0000000000000100;
assign   tb_i_aad[789]                        =   tb_i_aad[788];
assign   tb_i_rf_static_plaintext_length[789] =   64'h0000000000000280;
assign   tb_i_plaintext[789]                  =   tb_i_plaintext[788];
assign   tb_o_valid[789]                      =   1'b0;
assign   tb_o_sop[789]                        =   1'b0;
assign   tb_o_ciphertext[789]                 =   tb_o_ciphertext[788];
assign   tb_o_tag_ready[789]                  =   1'b0;
assign   tb_o_tag[789]                        =   tb_o_tag[788];

// CLK no. 790/1240
// *************************************************
assign   tb_i_valid[790]                      =   1'b0;
assign   tb_i_reset[790]                      =   1'b0;
assign   tb_i_sop[790]                        =   1'b0;
assign   tb_i_key_update[790]                 =   1'b0;
assign   tb_i_key[790]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[790]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[790]               =   1'b0;
assign   tb_i_rf_static_encrypt[790]          =   1'b1;
assign   tb_i_clear_fault_flags[790]          =   1'b0;
assign   tb_i_rf_static_aad_length[790]       =   64'h0000000000000100;
assign   tb_i_aad[790]                        =   tb_i_aad[789];
assign   tb_i_rf_static_plaintext_length[790] =   64'h0000000000000280;
assign   tb_i_plaintext[790]                  =   tb_i_plaintext[789];
assign   tb_o_valid[790]                      =   1'b0;
assign   tb_o_sop[790]                        =   1'b0;
assign   tb_o_ciphertext[790]                 =   tb_o_ciphertext[789];
assign   tb_o_tag_ready[790]                  =   1'b0;
assign   tb_o_tag[790]                        =   tb_o_tag[789];

// CLK no. 791/1240
// *************************************************
assign   tb_i_valid[791]                      =   1'b0;
assign   tb_i_reset[791]                      =   1'b0;
assign   tb_i_sop[791]                        =   1'b0;
assign   tb_i_key_update[791]                 =   1'b0;
assign   tb_i_key[791]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[791]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[791]               =   1'b0;
assign   tb_i_rf_static_encrypt[791]          =   1'b1;
assign   tb_i_clear_fault_flags[791]          =   1'b0;
assign   tb_i_rf_static_aad_length[791]       =   64'h0000000000000100;
assign   tb_i_aad[791]                        =   tb_i_aad[790];
assign   tb_i_rf_static_plaintext_length[791] =   64'h0000000000000280;
assign   tb_i_plaintext[791]                  =   tb_i_plaintext[790];
assign   tb_o_valid[791]                      =   1'b0;
assign   tb_o_sop[791]                        =   1'b0;
assign   tb_o_ciphertext[791]                 =   tb_o_ciphertext[790];
assign   tb_o_tag_ready[791]                  =   1'b0;
assign   tb_o_tag[791]                        =   tb_o_tag[790];

// CLK no. 792/1240
// *************************************************
assign   tb_i_valid[792]                      =   1'b0;
assign   tb_i_reset[792]                      =   1'b0;
assign   tb_i_sop[792]                        =   1'b0;
assign   tb_i_key_update[792]                 =   1'b0;
assign   tb_i_key[792]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[792]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[792]               =   1'b0;
assign   tb_i_rf_static_encrypt[792]          =   1'b1;
assign   tb_i_clear_fault_flags[792]          =   1'b0;
assign   tb_i_rf_static_aad_length[792]       =   64'h0000000000000100;
assign   tb_i_aad[792]                        =   tb_i_aad[791];
assign   tb_i_rf_static_plaintext_length[792] =   64'h0000000000000280;
assign   tb_i_plaintext[792]                  =   tb_i_plaintext[791];
assign   tb_o_valid[792]                      =   1'b0;
assign   tb_o_sop[792]                        =   1'b0;
assign   tb_o_ciphertext[792]                 =   tb_o_ciphertext[791];
assign   tb_o_tag_ready[792]                  =   1'b0;
assign   tb_o_tag[792]                        =   tb_o_tag[791];

// CLK no. 793/1240
// *************************************************
assign   tb_i_valid[793]                      =   1'b0;
assign   tb_i_reset[793]                      =   1'b0;
assign   tb_i_sop[793]                        =   1'b0;
assign   tb_i_key_update[793]                 =   1'b0;
assign   tb_i_key[793]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[793]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[793]               =   1'b0;
assign   tb_i_rf_static_encrypt[793]          =   1'b1;
assign   tb_i_clear_fault_flags[793]          =   1'b0;
assign   tb_i_rf_static_aad_length[793]       =   64'h0000000000000100;
assign   tb_i_aad[793]                        =   tb_i_aad[792];
assign   tb_i_rf_static_plaintext_length[793] =   64'h0000000000000280;
assign   tb_i_plaintext[793]                  =   tb_i_plaintext[792];
assign   tb_o_valid[793]                      =   1'b0;
assign   tb_o_sop[793]                        =   1'b0;
assign   tb_o_ciphertext[793]                 =   tb_o_ciphertext[792];
assign   tb_o_tag_ready[793]                  =   1'b0;
assign   tb_o_tag[793]                        =   tb_o_tag[792];

// CLK no. 794/1240
// *************************************************
assign   tb_i_valid[794]                      =   1'b0;
assign   tb_i_reset[794]                      =   1'b0;
assign   tb_i_sop[794]                        =   1'b0;
assign   tb_i_key_update[794]                 =   1'b0;
assign   tb_i_key[794]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[794]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[794]               =   1'b0;
assign   tb_i_rf_static_encrypt[794]          =   1'b1;
assign   tb_i_clear_fault_flags[794]          =   1'b0;
assign   tb_i_rf_static_aad_length[794]       =   64'h0000000000000100;
assign   tb_i_aad[794]                        =   tb_i_aad[793];
assign   tb_i_rf_static_plaintext_length[794] =   64'h0000000000000280;
assign   tb_i_plaintext[794]                  =   tb_i_plaintext[793];
assign   tb_o_valid[794]                      =   1'b0;
assign   tb_o_sop[794]                        =   1'b0;
assign   tb_o_ciphertext[794]                 =   tb_o_ciphertext[793];
assign   tb_o_tag_ready[794]                  =   1'b0;
assign   tb_o_tag[794]                        =   tb_o_tag[793];

// CLK no. 795/1240
// *************************************************
assign   tb_i_valid[795]                      =   1'b0;
assign   tb_i_reset[795]                      =   1'b0;
assign   tb_i_sop[795]                        =   1'b0;
assign   tb_i_key_update[795]                 =   1'b0;
assign   tb_i_key[795]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[795]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[795]               =   1'b0;
assign   tb_i_rf_static_encrypt[795]          =   1'b1;
assign   tb_i_clear_fault_flags[795]          =   1'b0;
assign   tb_i_rf_static_aad_length[795]       =   64'h0000000000000100;
assign   tb_i_aad[795]                        =   tb_i_aad[794];
assign   tb_i_rf_static_plaintext_length[795] =   64'h0000000000000280;
assign   tb_i_plaintext[795]                  =   tb_i_plaintext[794];
assign   tb_o_valid[795]                      =   1'b0;
assign   tb_o_sop[795]                        =   1'b0;
assign   tb_o_ciphertext[795]                 =   tb_o_ciphertext[794];
assign   tb_o_tag_ready[795]                  =   1'b0;
assign   tb_o_tag[795]                        =   tb_o_tag[794];

// CLK no. 796/1240
// *************************************************
assign   tb_i_valid[796]                      =   1'b0;
assign   tb_i_reset[796]                      =   1'b0;
assign   tb_i_sop[796]                        =   1'b0;
assign   tb_i_key_update[796]                 =   1'b0;
assign   tb_i_key[796]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[796]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[796]               =   1'b0;
assign   tb_i_rf_static_encrypt[796]          =   1'b1;
assign   tb_i_clear_fault_flags[796]          =   1'b0;
assign   tb_i_rf_static_aad_length[796]       =   64'h0000000000000100;
assign   tb_i_aad[796]                        =   tb_i_aad[795];
assign   tb_i_rf_static_plaintext_length[796] =   64'h0000000000000280;
assign   tb_i_plaintext[796]                  =   tb_i_plaintext[795];
assign   tb_o_valid[796]                      =   1'b0;
assign   tb_o_sop[796]                        =   1'b0;
assign   tb_o_ciphertext[796]                 =   tb_o_ciphertext[795];
assign   tb_o_tag_ready[796]                  =   1'b0;
assign   tb_o_tag[796]                        =   tb_o_tag[795];

// CLK no. 797/1240
// *************************************************
assign   tb_i_valid[797]                      =   1'b0;
assign   tb_i_reset[797]                      =   1'b0;
assign   tb_i_sop[797]                        =   1'b0;
assign   tb_i_key_update[797]                 =   1'b0;
assign   tb_i_key[797]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[797]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[797]               =   1'b0;
assign   tb_i_rf_static_encrypt[797]          =   1'b1;
assign   tb_i_clear_fault_flags[797]          =   1'b0;
assign   tb_i_rf_static_aad_length[797]       =   64'h0000000000000100;
assign   tb_i_aad[797]                        =   tb_i_aad[796];
assign   tb_i_rf_static_plaintext_length[797] =   64'h0000000000000280;
assign   tb_i_plaintext[797]                  =   tb_i_plaintext[796];
assign   tb_o_valid[797]                      =   1'b0;
assign   tb_o_sop[797]                        =   1'b0;
assign   tb_o_ciphertext[797]                 =   tb_o_ciphertext[796];
assign   tb_o_tag_ready[797]                  =   1'b0;
assign   tb_o_tag[797]                        =   tb_o_tag[796];

// CLK no. 798/1240
// *************************************************
assign   tb_i_valid[798]                      =   1'b0;
assign   tb_i_reset[798]                      =   1'b0;
assign   tb_i_sop[798]                        =   1'b0;
assign   tb_i_key_update[798]                 =   1'b0;
assign   tb_i_key[798]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[798]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[798]               =   1'b0;
assign   tb_i_rf_static_encrypt[798]          =   1'b1;
assign   tb_i_clear_fault_flags[798]          =   1'b0;
assign   tb_i_rf_static_aad_length[798]       =   64'h0000000000000100;
assign   tb_i_aad[798]                        =   tb_i_aad[797];
assign   tb_i_rf_static_plaintext_length[798] =   64'h0000000000000280;
assign   tb_i_plaintext[798]                  =   tb_i_plaintext[797];
assign   tb_o_valid[798]                      =   1'b0;
assign   tb_o_sop[798]                        =   1'b0;
assign   tb_o_ciphertext[798]                 =   tb_o_ciphertext[797];
assign   tb_o_tag_ready[798]                  =   1'b0;
assign   tb_o_tag[798]                        =   tb_o_tag[797];

// CLK no. 799/1240
// *************************************************
assign   tb_i_valid[799]                      =   1'b0;
assign   tb_i_reset[799]                      =   1'b0;
assign   tb_i_sop[799]                        =   1'b0;
assign   tb_i_key_update[799]                 =   1'b0;
assign   tb_i_key[799]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[799]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[799]               =   1'b0;
assign   tb_i_rf_static_encrypt[799]          =   1'b1;
assign   tb_i_clear_fault_flags[799]          =   1'b0;
assign   tb_i_rf_static_aad_length[799]       =   64'h0000000000000100;
assign   tb_i_aad[799]                        =   tb_i_aad[798];
assign   tb_i_rf_static_plaintext_length[799] =   64'h0000000000000280;
assign   tb_i_plaintext[799]                  =   tb_i_plaintext[798];
assign   tb_o_valid[799]                      =   1'b0;
assign   tb_o_sop[799]                        =   1'b0;
assign   tb_o_ciphertext[799]                 =   tb_o_ciphertext[798];
assign   tb_o_tag_ready[799]                  =   1'b0;
assign   tb_o_tag[799]                        =   tb_o_tag[798];

// CLK no. 800/1240
// *************************************************
assign   tb_i_valid[800]                      =   1'b0;
assign   tb_i_reset[800]                      =   1'b0;
assign   tb_i_sop[800]                        =   1'b0;
assign   tb_i_key_update[800]                 =   1'b0;
assign   tb_i_key[800]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[800]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[800]               =   1'b0;
assign   tb_i_rf_static_encrypt[800]          =   1'b1;
assign   tb_i_clear_fault_flags[800]          =   1'b0;
assign   tb_i_rf_static_aad_length[800]       =   64'h0000000000000100;
assign   tb_i_aad[800]                        =   tb_i_aad[799];
assign   tb_i_rf_static_plaintext_length[800] =   64'h0000000000000280;
assign   tb_i_plaintext[800]                  =   tb_i_plaintext[799];
assign   tb_o_valid[800]                      =   1'b0;
assign   tb_o_sop[800]                        =   1'b0;
assign   tb_o_ciphertext[800]                 =   tb_o_ciphertext[799];
assign   tb_o_tag_ready[800]                  =   1'b0;
assign   tb_o_tag[800]                        =   tb_o_tag[799];

// CLK no. 801/1240
// *************************************************
assign   tb_i_valid[801]                      =   1'b0;
assign   tb_i_reset[801]                      =   1'b0;
assign   tb_i_sop[801]                        =   1'b0;
assign   tb_i_key_update[801]                 =   1'b0;
assign   tb_i_key[801]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[801]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[801]               =   1'b0;
assign   tb_i_rf_static_encrypt[801]          =   1'b1;
assign   tb_i_clear_fault_flags[801]          =   1'b0;
assign   tb_i_rf_static_aad_length[801]       =   64'h0000000000000100;
assign   tb_i_aad[801]                        =   tb_i_aad[800];
assign   tb_i_rf_static_plaintext_length[801] =   64'h0000000000000280;
assign   tb_i_plaintext[801]                  =   tb_i_plaintext[800];
assign   tb_o_valid[801]                      =   1'b0;
assign   tb_o_sop[801]                        =   1'b0;
assign   tb_o_ciphertext[801]                 =   tb_o_ciphertext[800];
assign   tb_o_tag_ready[801]                  =   1'b0;
assign   tb_o_tag[801]                        =   tb_o_tag[800];

// CLK no. 802/1240
// *************************************************
assign   tb_i_valid[802]                      =   1'b0;
assign   tb_i_reset[802]                      =   1'b0;
assign   tb_i_sop[802]                        =   1'b0;
assign   tb_i_key_update[802]                 =   1'b0;
assign   tb_i_key[802]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[802]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[802]               =   1'b0;
assign   tb_i_rf_static_encrypt[802]          =   1'b1;
assign   tb_i_clear_fault_flags[802]          =   1'b0;
assign   tb_i_rf_static_aad_length[802]       =   64'h0000000000000100;
assign   tb_i_aad[802]                        =   tb_i_aad[801];
assign   tb_i_rf_static_plaintext_length[802] =   64'h0000000000000280;
assign   tb_i_plaintext[802]                  =   tb_i_plaintext[801];
assign   tb_o_valid[802]                      =   1'b0;
assign   tb_o_sop[802]                        =   1'b0;
assign   tb_o_ciphertext[802]                 =   tb_o_ciphertext[801];
assign   tb_o_tag_ready[802]                  =   1'b0;
assign   tb_o_tag[802]                        =   tb_o_tag[801];

// CLK no. 803/1240
// *************************************************
assign   tb_i_valid[803]                      =   1'b0;
assign   tb_i_reset[803]                      =   1'b0;
assign   tb_i_sop[803]                        =   1'b0;
assign   tb_i_key_update[803]                 =   1'b0;
assign   tb_i_key[803]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[803]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[803]               =   1'b0;
assign   tb_i_rf_static_encrypt[803]          =   1'b1;
assign   tb_i_clear_fault_flags[803]          =   1'b0;
assign   tb_i_rf_static_aad_length[803]       =   64'h0000000000000100;
assign   tb_i_aad[803]                        =   tb_i_aad[802];
assign   tb_i_rf_static_plaintext_length[803] =   64'h0000000000000280;
assign   tb_i_plaintext[803]                  =   tb_i_plaintext[802];
assign   tb_o_valid[803]                      =   1'b0;
assign   tb_o_sop[803]                        =   1'b0;
assign   tb_o_ciphertext[803]                 =   tb_o_ciphertext[802];
assign   tb_o_tag_ready[803]                  =   1'b0;
assign   tb_o_tag[803]                        =   tb_o_tag[802];

// CLK no. 804/1240
// *************************************************
assign   tb_i_valid[804]                      =   1'b0;
assign   tb_i_reset[804]                      =   1'b0;
assign   tb_i_sop[804]                        =   1'b0;
assign   tb_i_key_update[804]                 =   1'b0;
assign   tb_i_key[804]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[804]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[804]               =   1'b0;
assign   tb_i_rf_static_encrypt[804]          =   1'b1;
assign   tb_i_clear_fault_flags[804]          =   1'b0;
assign   tb_i_rf_static_aad_length[804]       =   64'h0000000000000100;
assign   tb_i_aad[804]                        =   tb_i_aad[803];
assign   tb_i_rf_static_plaintext_length[804] =   64'h0000000000000280;
assign   tb_i_plaintext[804]                  =   tb_i_plaintext[803];
assign   tb_o_valid[804]                      =   1'b0;
assign   tb_o_sop[804]                        =   1'b0;
assign   tb_o_ciphertext[804]                 =   tb_o_ciphertext[803];
assign   tb_o_tag_ready[804]                  =   1'b0;
assign   tb_o_tag[804]                        =   tb_o_tag[803];

// CLK no. 805/1240
// *************************************************
assign   tb_i_valid[805]                      =   1'b0;
assign   tb_i_reset[805]                      =   1'b0;
assign   tb_i_sop[805]                        =   1'b0;
assign   tb_i_key_update[805]                 =   1'b0;
assign   tb_i_key[805]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[805]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[805]               =   1'b0;
assign   tb_i_rf_static_encrypt[805]          =   1'b1;
assign   tb_i_clear_fault_flags[805]          =   1'b0;
assign   tb_i_rf_static_aad_length[805]       =   64'h0000000000000100;
assign   tb_i_aad[805]                        =   tb_i_aad[804];
assign   tb_i_rf_static_plaintext_length[805] =   64'h0000000000000280;
assign   tb_i_plaintext[805]                  =   tb_i_plaintext[804];
assign   tb_o_valid[805]                      =   1'b0;
assign   tb_o_sop[805]                        =   1'b0;
assign   tb_o_ciphertext[805]                 =   tb_o_ciphertext[804];
assign   tb_o_tag_ready[805]                  =   1'b0;
assign   tb_o_tag[805]                        =   tb_o_tag[804];

// CLK no. 806/1240
// *************************************************
assign   tb_i_valid[806]                      =   1'b0;
assign   tb_i_reset[806]                      =   1'b0;
assign   tb_i_sop[806]                        =   1'b0;
assign   tb_i_key_update[806]                 =   1'b0;
assign   tb_i_key[806]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[806]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[806]               =   1'b0;
assign   tb_i_rf_static_encrypt[806]          =   1'b1;
assign   tb_i_clear_fault_flags[806]          =   1'b0;
assign   tb_i_rf_static_aad_length[806]       =   64'h0000000000000100;
assign   tb_i_aad[806]                        =   tb_i_aad[805];
assign   tb_i_rf_static_plaintext_length[806] =   64'h0000000000000280;
assign   tb_i_plaintext[806]                  =   tb_i_plaintext[805];
assign   tb_o_valid[806]                      =   1'b0;
assign   tb_o_sop[806]                        =   1'b0;
assign   tb_o_ciphertext[806]                 =   tb_o_ciphertext[805];
assign   tb_o_tag_ready[806]                  =   1'b0;
assign   tb_o_tag[806]                        =   tb_o_tag[805];

// CLK no. 807/1240
// *************************************************
assign   tb_i_valid[807]                      =   1'b0;
assign   tb_i_reset[807]                      =   1'b0;
assign   tb_i_sop[807]                        =   1'b0;
assign   tb_i_key_update[807]                 =   1'b0;
assign   tb_i_key[807]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[807]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[807]               =   1'b0;
assign   tb_i_rf_static_encrypt[807]          =   1'b1;
assign   tb_i_clear_fault_flags[807]          =   1'b0;
assign   tb_i_rf_static_aad_length[807]       =   64'h0000000000000100;
assign   tb_i_aad[807]                        =   tb_i_aad[806];
assign   tb_i_rf_static_plaintext_length[807] =   64'h0000000000000280;
assign   tb_i_plaintext[807]                  =   tb_i_plaintext[806];
assign   tb_o_valid[807]                      =   1'b0;
assign   tb_o_sop[807]                        =   1'b0;
assign   tb_o_ciphertext[807]                 =   tb_o_ciphertext[806];
assign   tb_o_tag_ready[807]                  =   1'b0;
assign   tb_o_tag[807]                        =   tb_o_tag[806];

// CLK no. 808/1240
// *************************************************
assign   tb_i_valid[808]                      =   1'b0;
assign   tb_i_reset[808]                      =   1'b0;
assign   tb_i_sop[808]                        =   1'b0;
assign   tb_i_key_update[808]                 =   1'b0;
assign   tb_i_key[808]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[808]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[808]               =   1'b0;
assign   tb_i_rf_static_encrypt[808]          =   1'b1;
assign   tb_i_clear_fault_flags[808]          =   1'b0;
assign   tb_i_rf_static_aad_length[808]       =   64'h0000000000000100;
assign   tb_i_aad[808]                        =   tb_i_aad[807];
assign   tb_i_rf_static_plaintext_length[808] =   64'h0000000000000280;
assign   tb_i_plaintext[808]                  =   tb_i_plaintext[807];
assign   tb_o_valid[808]                      =   1'b0;
assign   tb_o_sop[808]                        =   1'b0;
assign   tb_o_ciphertext[808]                 =   tb_o_ciphertext[807];
assign   tb_o_tag_ready[808]                  =   1'b0;
assign   tb_o_tag[808]                        =   tb_o_tag[807];

// CLK no. 809/1240
// *************************************************
assign   tb_i_valid[809]                      =   1'b0;
assign   tb_i_reset[809]                      =   1'b0;
assign   tb_i_sop[809]                        =   1'b0;
assign   tb_i_key_update[809]                 =   1'b0;
assign   tb_i_key[809]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[809]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[809]               =   1'b0;
assign   tb_i_rf_static_encrypt[809]          =   1'b1;
assign   tb_i_clear_fault_flags[809]          =   1'b0;
assign   tb_i_rf_static_aad_length[809]       =   64'h0000000000000100;
assign   tb_i_aad[809]                        =   tb_i_aad[808];
assign   tb_i_rf_static_plaintext_length[809] =   64'h0000000000000280;
assign   tb_i_plaintext[809]                  =   tb_i_plaintext[808];
assign   tb_o_valid[809]                      =   1'b0;
assign   tb_o_sop[809]                        =   1'b0;
assign   tb_o_ciphertext[809]                 =   tb_o_ciphertext[808];
assign   tb_o_tag_ready[809]                  =   1'b0;
assign   tb_o_tag[809]                        =   tb_o_tag[808];

// CLK no. 810/1240
// *************************************************
assign   tb_i_valid[810]                      =   1'b0;
assign   tb_i_reset[810]                      =   1'b0;
assign   tb_i_sop[810]                        =   1'b0;
assign   tb_i_key_update[810]                 =   1'b0;
assign   tb_i_key[810]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[810]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[810]               =   1'b0;
assign   tb_i_rf_static_encrypt[810]          =   1'b1;
assign   tb_i_clear_fault_flags[810]          =   1'b0;
assign   tb_i_rf_static_aad_length[810]       =   64'h0000000000000100;
assign   tb_i_aad[810]                        =   tb_i_aad[809];
assign   tb_i_rf_static_plaintext_length[810] =   64'h0000000000000280;
assign   tb_i_plaintext[810]                  =   tb_i_plaintext[809];
assign   tb_o_valid[810]                      =   1'b0;
assign   tb_o_sop[810]                        =   1'b0;
assign   tb_o_ciphertext[810]                 =   tb_o_ciphertext[809];
assign   tb_o_tag_ready[810]                  =   1'b0;
assign   tb_o_tag[810]                        =   tb_o_tag[809];

// CLK no. 811/1240
// *************************************************
assign   tb_i_valid[811]                      =   1'b0;
assign   tb_i_reset[811]                      =   1'b0;
assign   tb_i_sop[811]                        =   1'b0;
assign   tb_i_key_update[811]                 =   1'b0;
assign   tb_i_key[811]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[811]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[811]               =   1'b0;
assign   tb_i_rf_static_encrypt[811]          =   1'b1;
assign   tb_i_clear_fault_flags[811]          =   1'b0;
assign   tb_i_rf_static_aad_length[811]       =   64'h0000000000000100;
assign   tb_i_aad[811]                        =   tb_i_aad[810];
assign   tb_i_rf_static_plaintext_length[811] =   64'h0000000000000280;
assign   tb_i_plaintext[811]                  =   tb_i_plaintext[810];
assign   tb_o_valid[811]                      =   1'b0;
assign   tb_o_sop[811]                        =   1'b0;
assign   tb_o_ciphertext[811]                 =   tb_o_ciphertext[810];
assign   tb_o_tag_ready[811]                  =   1'b0;
assign   tb_o_tag[811]                        =   tb_o_tag[810];

// CLK no. 812/1240
// *************************************************
assign   tb_i_valid[812]                      =   1'b0;
assign   tb_i_reset[812]                      =   1'b0;
assign   tb_i_sop[812]                        =   1'b0;
assign   tb_i_key_update[812]                 =   1'b0;
assign   tb_i_key[812]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[812]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[812]               =   1'b0;
assign   tb_i_rf_static_encrypt[812]          =   1'b1;
assign   tb_i_clear_fault_flags[812]          =   1'b0;
assign   tb_i_rf_static_aad_length[812]       =   64'h0000000000000100;
assign   tb_i_aad[812]                        =   tb_i_aad[811];
assign   tb_i_rf_static_plaintext_length[812] =   64'h0000000000000280;
assign   tb_i_plaintext[812]                  =   tb_i_plaintext[811];
assign   tb_o_valid[812]                      =   1'b0;
assign   tb_o_sop[812]                        =   1'b0;
assign   tb_o_ciphertext[812]                 =   tb_o_ciphertext[811];
assign   tb_o_tag_ready[812]                  =   1'b0;
assign   tb_o_tag[812]                        =   tb_o_tag[811];

// CLK no. 813/1240
// *************************************************
assign   tb_i_valid[813]                      =   1'b0;
assign   tb_i_reset[813]                      =   1'b0;
assign   tb_i_sop[813]                        =   1'b0;
assign   tb_i_key_update[813]                 =   1'b0;
assign   tb_i_key[813]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[813]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[813]               =   1'b0;
assign   tb_i_rf_static_encrypt[813]          =   1'b1;
assign   tb_i_clear_fault_flags[813]          =   1'b0;
assign   tb_i_rf_static_aad_length[813]       =   64'h0000000000000100;
assign   tb_i_aad[813]                        =   tb_i_aad[812];
assign   tb_i_rf_static_plaintext_length[813] =   64'h0000000000000280;
assign   tb_i_plaintext[813]                  =   tb_i_plaintext[812];
assign   tb_o_valid[813]                      =   1'b0;
assign   tb_o_sop[813]                        =   1'b0;
assign   tb_o_ciphertext[813]                 =   tb_o_ciphertext[812];
assign   tb_o_tag_ready[813]                  =   1'b0;
assign   tb_o_tag[813]                        =   tb_o_tag[812];

// CLK no. 814/1240
// *************************************************
assign   tb_i_valid[814]                      =   1'b0;
assign   tb_i_reset[814]                      =   1'b0;
assign   tb_i_sop[814]                        =   1'b0;
assign   tb_i_key_update[814]                 =   1'b0;
assign   tb_i_key[814]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[814]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[814]               =   1'b0;
assign   tb_i_rf_static_encrypt[814]          =   1'b1;
assign   tb_i_clear_fault_flags[814]          =   1'b0;
assign   tb_i_rf_static_aad_length[814]       =   64'h0000000000000100;
assign   tb_i_aad[814]                        =   tb_i_aad[813];
assign   tb_i_rf_static_plaintext_length[814] =   64'h0000000000000280;
assign   tb_i_plaintext[814]                  =   tb_i_plaintext[813];
assign   tb_o_valid[814]                      =   1'b1;
assign   tb_o_sop[814]                        =   1'b1;
assign   tb_o_ciphertext[814]                 =   256'h1c32bbe6f5bd85d6e7855baa99a0df3fcef5d89983e2e529a801a1ab42c1e9a0;
assign   tb_o_tag_ready[814]                  =   1'b0;
assign   tb_o_tag[814]                        =   tb_o_tag[813];

// CLK no. 815/1240
// *************************************************
assign   tb_i_valid[815]                      =   1'b0;
assign   tb_i_reset[815]                      =   1'b0;
assign   tb_i_sop[815]                        =   1'b0;
assign   tb_i_key_update[815]                 =   1'b0;
assign   tb_i_key[815]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[815]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[815]               =   1'b0;
assign   tb_i_rf_static_encrypt[815]          =   1'b1;
assign   tb_i_clear_fault_flags[815]          =   1'b0;
assign   tb_i_rf_static_aad_length[815]       =   64'h0000000000000100;
assign   tb_i_aad[815]                        =   tb_i_aad[814];
assign   tb_i_rf_static_plaintext_length[815] =   64'h0000000000000280;
assign   tb_i_plaintext[815]                  =   tb_i_plaintext[814];
assign   tb_o_valid[815]                      =   1'b1;
assign   tb_o_sop[815]                        =   1'b0;
assign   tb_o_ciphertext[815]                 =   256'h378f6c9856f726d20c1a43c1ce23f0fb4b97e29a9c4fd967cb2fdc4a6af7d44f;
assign   tb_o_tag_ready[815]                  =   1'b0;
assign   tb_o_tag[815]                        =   tb_o_tag[814];

// CLK no. 816/1240
// *************************************************
assign   tb_i_valid[816]                      =   1'b0;
assign   tb_i_reset[816]                      =   1'b0;
assign   tb_i_sop[816]                        =   1'b0;
assign   tb_i_key_update[816]                 =   1'b0;
assign   tb_i_key[816]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[816]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[816]               =   1'b0;
assign   tb_i_rf_static_encrypt[816]          =   1'b1;
assign   tb_i_clear_fault_flags[816]          =   1'b0;
assign   tb_i_rf_static_aad_length[816]       =   64'h0000000000000100;
assign   tb_i_aad[816]                        =   tb_i_aad[815];
assign   tb_i_rf_static_plaintext_length[816] =   64'h0000000000000280;
assign   tb_i_plaintext[816]                  =   tb_i_plaintext[815];
assign   tb_o_valid[816]                      =   1'b1;
assign   tb_o_sop[816]                        =   1'b0;
assign   tb_o_ciphertext[816]                 =   256'h84c2467e8ef7c5f19f6fb60954e4cd1d;
assign   tb_o_tag_ready[816]                  =   1'b0;
assign   tb_o_tag[816]                        =   tb_o_tag[815];

// CLK no. 817/1240
// *************************************************
assign   tb_i_valid[817]                      =   1'b0;
assign   tb_i_reset[817]                      =   1'b0;
assign   tb_i_sop[817]                        =   1'b0;
assign   tb_i_key_update[817]                 =   1'b0;
assign   tb_i_key[817]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[817]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[817]               =   1'b0;
assign   tb_i_rf_static_encrypt[817]          =   1'b1;
assign   tb_i_clear_fault_flags[817]          =   1'b0;
assign   tb_i_rf_static_aad_length[817]       =   64'h0000000000000100;
assign   tb_i_aad[817]                        =   tb_i_aad[816];
assign   tb_i_rf_static_plaintext_length[817] =   64'h0000000000000280;
assign   tb_i_plaintext[817]                  =   tb_i_plaintext[816];
assign   tb_o_valid[817]                      =   1'b0;
assign   tb_o_sop[817]                        =   1'b0;
assign   tb_o_ciphertext[817]                 =   tb_o_ciphertext[816];
assign   tb_o_tag_ready[817]                  =   1'b0;
assign   tb_o_tag[817]                        =   tb_o_tag[816];

// CLK no. 818/1240
// *************************************************
assign   tb_i_valid[818]                      =   1'b0;
assign   tb_i_reset[818]                      =   1'b0;
assign   tb_i_sop[818]                        =   1'b0;
assign   tb_i_key_update[818]                 =   1'b0;
assign   tb_i_key[818]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[818]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[818]               =   1'b0;
assign   tb_i_rf_static_encrypt[818]          =   1'b1;
assign   tb_i_clear_fault_flags[818]          =   1'b0;
assign   tb_i_rf_static_aad_length[818]       =   64'h0000000000000100;
assign   tb_i_aad[818]                        =   tb_i_aad[817];
assign   tb_i_rf_static_plaintext_length[818] =   64'h0000000000000280;
assign   tb_i_plaintext[818]                  =   tb_i_plaintext[817];
assign   tb_o_valid[818]                      =   1'b0;
assign   tb_o_sop[818]                        =   1'b0;
assign   tb_o_ciphertext[818]                 =   tb_o_ciphertext[817];
assign   tb_o_tag_ready[818]                  =   1'b0;
assign   tb_o_tag[818]                        =   tb_o_tag[817];

// CLK no. 819/1240
// *************************************************
assign   tb_i_valid[819]                      =   1'b0;
assign   tb_i_reset[819]                      =   1'b0;
assign   tb_i_sop[819]                        =   1'b0;
assign   tb_i_key_update[819]                 =   1'b0;
assign   tb_i_key[819]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[819]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[819]               =   1'b0;
assign   tb_i_rf_static_encrypt[819]          =   1'b1;
assign   tb_i_clear_fault_flags[819]          =   1'b0;
assign   tb_i_rf_static_aad_length[819]       =   64'h0000000000000100;
assign   tb_i_aad[819]                        =   tb_i_aad[818];
assign   tb_i_rf_static_plaintext_length[819] =   64'h0000000000000280;
assign   tb_i_plaintext[819]                  =   tb_i_plaintext[818];
assign   tb_o_valid[819]                      =   1'b0;
assign   tb_o_sop[819]                        =   1'b0;
assign   tb_o_ciphertext[819]                 =   tb_o_ciphertext[818];
assign   tb_o_tag_ready[819]                  =   1'b0;
assign   tb_o_tag[819]                        =   tb_o_tag[818];

// CLK no. 820/1240
// *************************************************
assign   tb_i_valid[820]                      =   1'b0;
assign   tb_i_reset[820]                      =   1'b0;
assign   tb_i_sop[820]                        =   1'b0;
assign   tb_i_key_update[820]                 =   1'b0;
assign   tb_i_key[820]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[820]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[820]               =   1'b0;
assign   tb_i_rf_static_encrypt[820]          =   1'b1;
assign   tb_i_clear_fault_flags[820]          =   1'b0;
assign   tb_i_rf_static_aad_length[820]       =   64'h0000000000000100;
assign   tb_i_aad[820]                        =   tb_i_aad[819];
assign   tb_i_rf_static_plaintext_length[820] =   64'h0000000000000280;
assign   tb_i_plaintext[820]                  =   tb_i_plaintext[819];
assign   tb_o_valid[820]                      =   1'b0;
assign   tb_o_sop[820]                        =   1'b0;
assign   tb_o_ciphertext[820]                 =   tb_o_ciphertext[819];
assign   tb_o_tag_ready[820]                  =   1'b0;
assign   tb_o_tag[820]                        =   tb_o_tag[819];

// CLK no. 821/1240
// *************************************************
assign   tb_i_valid[821]                      =   1'b0;
assign   tb_i_reset[821]                      =   1'b0;
assign   tb_i_sop[821]                        =   1'b0;
assign   tb_i_key_update[821]                 =   1'b0;
assign   tb_i_key[821]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[821]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[821]               =   1'b0;
assign   tb_i_rf_static_encrypt[821]          =   1'b1;
assign   tb_i_clear_fault_flags[821]          =   1'b0;
assign   tb_i_rf_static_aad_length[821]       =   64'h0000000000000100;
assign   tb_i_aad[821]                        =   tb_i_aad[820];
assign   tb_i_rf_static_plaintext_length[821] =   64'h0000000000000280;
assign   tb_i_plaintext[821]                  =   tb_i_plaintext[820];
assign   tb_o_valid[821]                      =   1'b0;
assign   tb_o_sop[821]                        =   1'b0;
assign   tb_o_ciphertext[821]                 =   tb_o_ciphertext[820];
assign   tb_o_tag_ready[821]                  =   1'b0;
assign   tb_o_tag[821]                        =   tb_o_tag[820];

// CLK no. 822/1240
// *************************************************
assign   tb_i_valid[822]                      =   1'b0;
assign   tb_i_reset[822]                      =   1'b0;
assign   tb_i_sop[822]                        =   1'b0;
assign   tb_i_key_update[822]                 =   1'b0;
assign   tb_i_key[822]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[822]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[822]               =   1'b0;
assign   tb_i_rf_static_encrypt[822]          =   1'b1;
assign   tb_i_clear_fault_flags[822]          =   1'b0;
assign   tb_i_rf_static_aad_length[822]       =   64'h0000000000000100;
assign   tb_i_aad[822]                        =   tb_i_aad[821];
assign   tb_i_rf_static_plaintext_length[822] =   64'h0000000000000280;
assign   tb_i_plaintext[822]                  =   tb_i_plaintext[821];
assign   tb_o_valid[822]                      =   1'b0;
assign   tb_o_sop[822]                        =   1'b0;
assign   tb_o_ciphertext[822]                 =   tb_o_ciphertext[821];
assign   tb_o_tag_ready[822]                  =   1'b0;
assign   tb_o_tag[822]                        =   tb_o_tag[821];

// CLK no. 823/1240
// *************************************************
assign   tb_i_valid[823]                      =   1'b0;
assign   tb_i_reset[823]                      =   1'b0;
assign   tb_i_sop[823]                        =   1'b0;
assign   tb_i_key_update[823]                 =   1'b0;
assign   tb_i_key[823]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[823]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[823]               =   1'b0;
assign   tb_i_rf_static_encrypt[823]          =   1'b1;
assign   tb_i_clear_fault_flags[823]          =   1'b0;
assign   tb_i_rf_static_aad_length[823]       =   64'h0000000000000100;
assign   tb_i_aad[823]                        =   tb_i_aad[822];
assign   tb_i_rf_static_plaintext_length[823] =   64'h0000000000000280;
assign   tb_i_plaintext[823]                  =   tb_i_plaintext[822];
assign   tb_o_valid[823]                      =   1'b0;
assign   tb_o_sop[823]                        =   1'b0;
assign   tb_o_ciphertext[823]                 =   tb_o_ciphertext[822];
assign   tb_o_tag_ready[823]                  =   1'b0;
assign   tb_o_tag[823]                        =   tb_o_tag[822];

// CLK no. 824/1240
// *************************************************
assign   tb_i_valid[824]                      =   1'b0;
assign   tb_i_reset[824]                      =   1'b0;
assign   tb_i_sop[824]                        =   1'b0;
assign   tb_i_key_update[824]                 =   1'b0;
assign   tb_i_key[824]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[824]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[824]               =   1'b0;
assign   tb_i_rf_static_encrypt[824]          =   1'b1;
assign   tb_i_clear_fault_flags[824]          =   1'b0;
assign   tb_i_rf_static_aad_length[824]       =   64'h0000000000000100;
assign   tb_i_aad[824]                        =   tb_i_aad[823];
assign   tb_i_rf_static_plaintext_length[824] =   64'h0000000000000280;
assign   tb_i_plaintext[824]                  =   tb_i_plaintext[823];
assign   tb_o_valid[824]                      =   1'b0;
assign   tb_o_sop[824]                        =   1'b0;
assign   tb_o_ciphertext[824]                 =   tb_o_ciphertext[823];
assign   tb_o_tag_ready[824]                  =   1'b1;
assign   tb_o_tag[824]                        =   128'hdf08365eba6c9f7e028ad3ac9e427a55;

// CLK no. 825/1240
// *************************************************
assign   tb_i_valid[825]                      =   1'b0;
assign   tb_i_reset[825]                      =   1'b0;
assign   tb_i_sop[825]                        =   1'b0;
assign   tb_i_key_update[825]                 =   1'b0;
assign   tb_i_key[825]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[825]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[825]               =   1'b0;
assign   tb_i_rf_static_encrypt[825]          =   1'b1;
assign   tb_i_clear_fault_flags[825]          =   1'b0;
assign   tb_i_rf_static_aad_length[825]       =   64'h0000000000000100;
assign   tb_i_aad[825]                        =   tb_i_aad[824];
assign   tb_i_rf_static_plaintext_length[825] =   64'h0000000000000280;
assign   tb_i_plaintext[825]                  =   tb_i_plaintext[824];
assign   tb_o_valid[825]                      =   1'b0;
assign   tb_o_sop[825]                        =   1'b0;
assign   tb_o_ciphertext[825]                 =   tb_o_ciphertext[824];
assign   tb_o_tag_ready[825]                  =   1'b0;
assign   tb_o_tag[825]                        =   tb_o_tag[824];

// CLK no. 826/1240
// *************************************************
assign   tb_i_valid[826]                      =   1'b0;
assign   tb_i_reset[826]                      =   1'b0;
assign   tb_i_sop[826]                        =   1'b0;
assign   tb_i_key_update[826]                 =   1'b0;
assign   tb_i_key[826]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[826]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[826]               =   1'b0;
assign   tb_i_rf_static_encrypt[826]          =   1'b1;
assign   tb_i_clear_fault_flags[826]          =   1'b0;
assign   tb_i_rf_static_aad_length[826]       =   64'h0000000000000100;
assign   tb_i_aad[826]                        =   tb_i_aad[825];
assign   tb_i_rf_static_plaintext_length[826] =   64'h0000000000000280;
assign   tb_i_plaintext[826]                  =   tb_i_plaintext[825];
assign   tb_o_valid[826]                      =   1'b0;
assign   tb_o_sop[826]                        =   1'b0;
assign   tb_o_ciphertext[826]                 =   tb_o_ciphertext[825];
assign   tb_o_tag_ready[826]                  =   1'b0;
assign   tb_o_tag[826]                        =   tb_o_tag[825];

// CLK no. 827/1240
// *************************************************
assign   tb_i_valid[827]                      =   1'b0;
assign   tb_i_reset[827]                      =   1'b0;
assign   tb_i_sop[827]                        =   1'b1;
assign   tb_i_key_update[827]                 =   1'b0;
assign   tb_i_key[827]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[827]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[827]               =   1'b0;
assign   tb_i_rf_static_encrypt[827]          =   1'b1;
assign   tb_i_clear_fault_flags[827]          =   1'b0;
assign   tb_i_rf_static_aad_length[827]       =   64'h0000000000000100;
assign   tb_i_aad[827]                        =   tb_i_aad[826];
assign   tb_i_rf_static_plaintext_length[827] =   64'h0000000000000280;
assign   tb_i_plaintext[827]                  =   tb_i_plaintext[826];
assign   tb_o_valid[827]                      =   1'b0;
assign   tb_o_sop[827]                        =   1'b0;
assign   tb_o_ciphertext[827]                 =   tb_o_ciphertext[826];
assign   tb_o_tag_ready[827]                  =   1'b0;
assign   tb_o_tag[827]                        =   tb_o_tag[826];

// CLK no. 828/1240
// *************************************************
assign   tb_i_valid[828]                      =   1'b1;
assign   tb_i_reset[828]                      =   1'b0;
assign   tb_i_sop[828]                        =   1'b0;
assign   tb_i_key_update[828]                 =   1'b0;
assign   tb_i_key[828]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[828]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[828]               =   1'b0;
assign   tb_i_rf_static_encrypt[828]          =   1'b1;
assign   tb_i_clear_fault_flags[828]          =   1'b0;
assign   tb_i_rf_static_aad_length[828]       =   64'h0000000000000100;
assign   tb_i_aad[828]                        =   256'h947006894d6bd005bc04cc226ec044ab27349eb65c46469d870a8e1f67258092;
assign   tb_i_rf_static_plaintext_length[828] =   64'h0000000000000280;
assign   tb_i_plaintext[828]                  =   tb_i_plaintext[827];
assign   tb_o_valid[828]                      =   1'b0;
assign   tb_o_sop[828]                        =   1'b0;
assign   tb_o_ciphertext[828]                 =   tb_o_ciphertext[827];
assign   tb_o_tag_ready[828]                  =   1'b0;
assign   tb_o_tag[828]                        =   tb_o_tag[827];

// CLK no. 829/1240
// *************************************************
assign   tb_i_valid[829]                      =   1'b1;
assign   tb_i_reset[829]                      =   1'b0;
assign   tb_i_sop[829]                        =   1'b0;
assign   tb_i_key_update[829]                 =   1'b0;
assign   tb_i_key[829]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[829]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[829]               =   1'b0;
assign   tb_i_rf_static_encrypt[829]          =   1'b1;
assign   tb_i_clear_fault_flags[829]          =   1'b0;
assign   tb_i_rf_static_aad_length[829]       =   64'h0000000000000100;
assign   tb_i_aad[829]                        =   tb_i_aad[828];
assign   tb_i_rf_static_plaintext_length[829] =   64'h0000000000000280;
assign   tb_i_plaintext[829]                  =   256'h797f90e70c85a2361a7cb8954faaae102f215f6b973dcf07c7cd9a01b62438e8;
assign   tb_o_valid[829]                      =   1'b0;
assign   tb_o_sop[829]                        =   1'b0;
assign   tb_o_ciphertext[829]                 =   tb_o_ciphertext[828];
assign   tb_o_tag_ready[829]                  =   1'b0;
assign   tb_o_tag[829]                        =   tb_o_tag[828];

// CLK no. 830/1240
// *************************************************
assign   tb_i_valid[830]                      =   1'b1;
assign   tb_i_reset[830]                      =   1'b0;
assign   tb_i_sop[830]                        =   1'b0;
assign   tb_i_key_update[830]                 =   1'b0;
assign   tb_i_key[830]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[830]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[830]               =   1'b0;
assign   tb_i_rf_static_encrypt[830]          =   1'b1;
assign   tb_i_clear_fault_flags[830]          =   1'b0;
assign   tb_i_rf_static_aad_length[830]       =   64'h0000000000000100;
assign   tb_i_aad[830]                        =   tb_i_aad[829];
assign   tb_i_rf_static_plaintext_length[830] =   64'h0000000000000280;
assign   tb_i_plaintext[830]                  =   256'h894f15134bd6c98cf1460103479aa13c5b63b365c8e31825062b6e7ec0fe82db;
assign   tb_o_valid[830]                      =   1'b0;
assign   tb_o_sop[830]                        =   1'b0;
assign   tb_o_ciphertext[830]                 =   tb_o_ciphertext[829];
assign   tb_o_tag_ready[830]                  =   1'b0;
assign   tb_o_tag[830]                        =   tb_o_tag[829];

// CLK no. 831/1240
// *************************************************
assign   tb_i_valid[831]                      =   1'b1;
assign   tb_i_reset[831]                      =   1'b0;
assign   tb_i_sop[831]                        =   1'b0;
assign   tb_i_key_update[831]                 =   1'b0;
assign   tb_i_key[831]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[831]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[831]               =   1'b0;
assign   tb_i_rf_static_encrypt[831]          =   1'b1;
assign   tb_i_clear_fault_flags[831]          =   1'b0;
assign   tb_i_rf_static_aad_length[831]       =   64'h0000000000000100;
assign   tb_i_aad[831]                        =   tb_i_aad[830];
assign   tb_i_rf_static_plaintext_length[831] =   64'h0000000000000280;
assign   tb_i_plaintext[831]                  =   256'h8487857d9be77646aabd912921ec0513;
assign   tb_o_valid[831]                      =   1'b0;
assign   tb_o_sop[831]                        =   1'b0;
assign   tb_o_ciphertext[831]                 =   tb_o_ciphertext[830];
assign   tb_o_tag_ready[831]                  =   1'b0;
assign   tb_o_tag[831]                        =   tb_o_tag[830];

// CLK no. 832/1240
// *************************************************
assign   tb_i_valid[832]                      =   1'b0;
assign   tb_i_reset[832]                      =   1'b0;
assign   tb_i_sop[832]                        =   1'b0;
assign   tb_i_key_update[832]                 =   1'b0;
assign   tb_i_key[832]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[832]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[832]               =   1'b0;
assign   tb_i_rf_static_encrypt[832]          =   1'b1;
assign   tb_i_clear_fault_flags[832]          =   1'b0;
assign   tb_i_rf_static_aad_length[832]       =   64'h0000000000000100;
assign   tb_i_aad[832]                        =   tb_i_aad[831];
assign   tb_i_rf_static_plaintext_length[832] =   64'h0000000000000280;
assign   tb_i_plaintext[832]                  =   tb_i_plaintext[831];
assign   tb_o_valid[832]                      =   1'b0;
assign   tb_o_sop[832]                        =   1'b0;
assign   tb_o_ciphertext[832]                 =   tb_o_ciphertext[831];
assign   tb_o_tag_ready[832]                  =   1'b0;
assign   tb_o_tag[832]                        =   tb_o_tag[831];

// CLK no. 833/1240
// *************************************************
assign   tb_i_valid[833]                      =   1'b0;
assign   tb_i_reset[833]                      =   1'b0;
assign   tb_i_sop[833]                        =   1'b0;
assign   tb_i_key_update[833]                 =   1'b0;
assign   tb_i_key[833]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[833]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[833]               =   1'b0;
assign   tb_i_rf_static_encrypt[833]          =   1'b1;
assign   tb_i_clear_fault_flags[833]          =   1'b0;
assign   tb_i_rf_static_aad_length[833]       =   64'h0000000000000100;
assign   tb_i_aad[833]                        =   tb_i_aad[832];
assign   tb_i_rf_static_plaintext_length[833] =   64'h0000000000000280;
assign   tb_i_plaintext[833]                  =   tb_i_plaintext[832];
assign   tb_o_valid[833]                      =   1'b0;
assign   tb_o_sop[833]                        =   1'b0;
assign   tb_o_ciphertext[833]                 =   tb_o_ciphertext[832];
assign   tb_o_tag_ready[833]                  =   1'b0;
assign   tb_o_tag[833]                        =   tb_o_tag[832];

// CLK no. 834/1240
// *************************************************
assign   tb_i_valid[834]                      =   1'b0;
assign   tb_i_reset[834]                      =   1'b0;
assign   tb_i_sop[834]                        =   1'b0;
assign   tb_i_key_update[834]                 =   1'b0;
assign   tb_i_key[834]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[834]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[834]               =   1'b0;
assign   tb_i_rf_static_encrypt[834]          =   1'b1;
assign   tb_i_clear_fault_flags[834]          =   1'b0;
assign   tb_i_rf_static_aad_length[834]       =   64'h0000000000000100;
assign   tb_i_aad[834]                        =   tb_i_aad[833];
assign   tb_i_rf_static_plaintext_length[834] =   64'h0000000000000280;
assign   tb_i_plaintext[834]                  =   tb_i_plaintext[833];
assign   tb_o_valid[834]                      =   1'b0;
assign   tb_o_sop[834]                        =   1'b0;
assign   tb_o_ciphertext[834]                 =   tb_o_ciphertext[833];
assign   tb_o_tag_ready[834]                  =   1'b0;
assign   tb_o_tag[834]                        =   tb_o_tag[833];

// CLK no. 835/1240
// *************************************************
assign   tb_i_valid[835]                      =   1'b0;
assign   tb_i_reset[835]                      =   1'b0;
assign   tb_i_sop[835]                        =   1'b0;
assign   tb_i_key_update[835]                 =   1'b0;
assign   tb_i_key[835]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[835]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[835]               =   1'b0;
assign   tb_i_rf_static_encrypt[835]          =   1'b1;
assign   tb_i_clear_fault_flags[835]          =   1'b0;
assign   tb_i_rf_static_aad_length[835]       =   64'h0000000000000100;
assign   tb_i_aad[835]                        =   tb_i_aad[834];
assign   tb_i_rf_static_plaintext_length[835] =   64'h0000000000000280;
assign   tb_i_plaintext[835]                  =   tb_i_plaintext[834];
assign   tb_o_valid[835]                      =   1'b0;
assign   tb_o_sop[835]                        =   1'b0;
assign   tb_o_ciphertext[835]                 =   tb_o_ciphertext[834];
assign   tb_o_tag_ready[835]                  =   1'b0;
assign   tb_o_tag[835]                        =   tb_o_tag[834];

// CLK no. 836/1240
// *************************************************
assign   tb_i_valid[836]                      =   1'b0;
assign   tb_i_reset[836]                      =   1'b0;
assign   tb_i_sop[836]                        =   1'b0;
assign   tb_i_key_update[836]                 =   1'b0;
assign   tb_i_key[836]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[836]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[836]               =   1'b0;
assign   tb_i_rf_static_encrypt[836]          =   1'b1;
assign   tb_i_clear_fault_flags[836]          =   1'b0;
assign   tb_i_rf_static_aad_length[836]       =   64'h0000000000000100;
assign   tb_i_aad[836]                        =   tb_i_aad[835];
assign   tb_i_rf_static_plaintext_length[836] =   64'h0000000000000280;
assign   tb_i_plaintext[836]                  =   tb_i_plaintext[835];
assign   tb_o_valid[836]                      =   1'b0;
assign   tb_o_sop[836]                        =   1'b0;
assign   tb_o_ciphertext[836]                 =   tb_o_ciphertext[835];
assign   tb_o_tag_ready[836]                  =   1'b0;
assign   tb_o_tag[836]                        =   tb_o_tag[835];

// CLK no. 837/1240
// *************************************************
assign   tb_i_valid[837]                      =   1'b0;
assign   tb_i_reset[837]                      =   1'b0;
assign   tb_i_sop[837]                        =   1'b0;
assign   tb_i_key_update[837]                 =   1'b0;
assign   tb_i_key[837]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[837]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[837]               =   1'b0;
assign   tb_i_rf_static_encrypt[837]          =   1'b1;
assign   tb_i_clear_fault_flags[837]          =   1'b0;
assign   tb_i_rf_static_aad_length[837]       =   64'h0000000000000100;
assign   tb_i_aad[837]                        =   tb_i_aad[836];
assign   tb_i_rf_static_plaintext_length[837] =   64'h0000000000000280;
assign   tb_i_plaintext[837]                  =   tb_i_plaintext[836];
assign   tb_o_valid[837]                      =   1'b0;
assign   tb_o_sop[837]                        =   1'b0;
assign   tb_o_ciphertext[837]                 =   tb_o_ciphertext[836];
assign   tb_o_tag_ready[837]                  =   1'b0;
assign   tb_o_tag[837]                        =   tb_o_tag[836];

// CLK no. 838/1240
// *************************************************
assign   tb_i_valid[838]                      =   1'b0;
assign   tb_i_reset[838]                      =   1'b0;
assign   tb_i_sop[838]                        =   1'b0;
assign   tb_i_key_update[838]                 =   1'b0;
assign   tb_i_key[838]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[838]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[838]               =   1'b0;
assign   tb_i_rf_static_encrypt[838]          =   1'b1;
assign   tb_i_clear_fault_flags[838]          =   1'b0;
assign   tb_i_rf_static_aad_length[838]       =   64'h0000000000000100;
assign   tb_i_aad[838]                        =   tb_i_aad[837];
assign   tb_i_rf_static_plaintext_length[838] =   64'h0000000000000280;
assign   tb_i_plaintext[838]                  =   tb_i_plaintext[837];
assign   tb_o_valid[838]                      =   1'b0;
assign   tb_o_sop[838]                        =   1'b0;
assign   tb_o_ciphertext[838]                 =   tb_o_ciphertext[837];
assign   tb_o_tag_ready[838]                  =   1'b0;
assign   tb_o_tag[838]                        =   tb_o_tag[837];

// CLK no. 839/1240
// *************************************************
assign   tb_i_valid[839]                      =   1'b0;
assign   tb_i_reset[839]                      =   1'b0;
assign   tb_i_sop[839]                        =   1'b0;
assign   tb_i_key_update[839]                 =   1'b0;
assign   tb_i_key[839]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[839]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[839]               =   1'b0;
assign   tb_i_rf_static_encrypt[839]          =   1'b1;
assign   tb_i_clear_fault_flags[839]          =   1'b0;
assign   tb_i_rf_static_aad_length[839]       =   64'h0000000000000100;
assign   tb_i_aad[839]                        =   tb_i_aad[838];
assign   tb_i_rf_static_plaintext_length[839] =   64'h0000000000000280;
assign   tb_i_plaintext[839]                  =   tb_i_plaintext[838];
assign   tb_o_valid[839]                      =   1'b0;
assign   tb_o_sop[839]                        =   1'b0;
assign   tb_o_ciphertext[839]                 =   tb_o_ciphertext[838];
assign   tb_o_tag_ready[839]                  =   1'b0;
assign   tb_o_tag[839]                        =   tb_o_tag[838];

// CLK no. 840/1240
// *************************************************
assign   tb_i_valid[840]                      =   1'b0;
assign   tb_i_reset[840]                      =   1'b0;
assign   tb_i_sop[840]                        =   1'b0;
assign   tb_i_key_update[840]                 =   1'b0;
assign   tb_i_key[840]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[840]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[840]               =   1'b0;
assign   tb_i_rf_static_encrypt[840]          =   1'b1;
assign   tb_i_clear_fault_flags[840]          =   1'b0;
assign   tb_i_rf_static_aad_length[840]       =   64'h0000000000000100;
assign   tb_i_aad[840]                        =   tb_i_aad[839];
assign   tb_i_rf_static_plaintext_length[840] =   64'h0000000000000280;
assign   tb_i_plaintext[840]                  =   tb_i_plaintext[839];
assign   tb_o_valid[840]                      =   1'b0;
assign   tb_o_sop[840]                        =   1'b0;
assign   tb_o_ciphertext[840]                 =   tb_o_ciphertext[839];
assign   tb_o_tag_ready[840]                  =   1'b0;
assign   tb_o_tag[840]                        =   tb_o_tag[839];

// CLK no. 841/1240
// *************************************************
assign   tb_i_valid[841]                      =   1'b0;
assign   tb_i_reset[841]                      =   1'b0;
assign   tb_i_sop[841]                        =   1'b0;
assign   tb_i_key_update[841]                 =   1'b0;
assign   tb_i_key[841]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[841]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[841]               =   1'b0;
assign   tb_i_rf_static_encrypt[841]          =   1'b1;
assign   tb_i_clear_fault_flags[841]          =   1'b0;
assign   tb_i_rf_static_aad_length[841]       =   64'h0000000000000100;
assign   tb_i_aad[841]                        =   tb_i_aad[840];
assign   tb_i_rf_static_plaintext_length[841] =   64'h0000000000000280;
assign   tb_i_plaintext[841]                  =   tb_i_plaintext[840];
assign   tb_o_valid[841]                      =   1'b0;
assign   tb_o_sop[841]                        =   1'b0;
assign   tb_o_ciphertext[841]                 =   tb_o_ciphertext[840];
assign   tb_o_tag_ready[841]                  =   1'b0;
assign   tb_o_tag[841]                        =   tb_o_tag[840];

// CLK no. 842/1240
// *************************************************
assign   tb_i_valid[842]                      =   1'b0;
assign   tb_i_reset[842]                      =   1'b0;
assign   tb_i_sop[842]                        =   1'b0;
assign   tb_i_key_update[842]                 =   1'b0;
assign   tb_i_key[842]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[842]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[842]               =   1'b0;
assign   tb_i_rf_static_encrypt[842]          =   1'b1;
assign   tb_i_clear_fault_flags[842]          =   1'b0;
assign   tb_i_rf_static_aad_length[842]       =   64'h0000000000000100;
assign   tb_i_aad[842]                        =   tb_i_aad[841];
assign   tb_i_rf_static_plaintext_length[842] =   64'h0000000000000280;
assign   tb_i_plaintext[842]                  =   tb_i_plaintext[841];
assign   tb_o_valid[842]                      =   1'b0;
assign   tb_o_sop[842]                        =   1'b0;
assign   tb_o_ciphertext[842]                 =   tb_o_ciphertext[841];
assign   tb_o_tag_ready[842]                  =   1'b0;
assign   tb_o_tag[842]                        =   tb_o_tag[841];

// CLK no. 843/1240
// *************************************************
assign   tb_i_valid[843]                      =   1'b0;
assign   tb_i_reset[843]                      =   1'b0;
assign   tb_i_sop[843]                        =   1'b0;
assign   tb_i_key_update[843]                 =   1'b0;
assign   tb_i_key[843]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[843]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[843]               =   1'b0;
assign   tb_i_rf_static_encrypt[843]          =   1'b1;
assign   tb_i_clear_fault_flags[843]          =   1'b0;
assign   tb_i_rf_static_aad_length[843]       =   64'h0000000000000100;
assign   tb_i_aad[843]                        =   tb_i_aad[842];
assign   tb_i_rf_static_plaintext_length[843] =   64'h0000000000000280;
assign   tb_i_plaintext[843]                  =   tb_i_plaintext[842];
assign   tb_o_valid[843]                      =   1'b0;
assign   tb_o_sop[843]                        =   1'b0;
assign   tb_o_ciphertext[843]                 =   tb_o_ciphertext[842];
assign   tb_o_tag_ready[843]                  =   1'b0;
assign   tb_o_tag[843]                        =   tb_o_tag[842];

// CLK no. 844/1240
// *************************************************
assign   tb_i_valid[844]                      =   1'b0;
assign   tb_i_reset[844]                      =   1'b0;
assign   tb_i_sop[844]                        =   1'b0;
assign   tb_i_key_update[844]                 =   1'b0;
assign   tb_i_key[844]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[844]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[844]               =   1'b0;
assign   tb_i_rf_static_encrypt[844]          =   1'b1;
assign   tb_i_clear_fault_flags[844]          =   1'b0;
assign   tb_i_rf_static_aad_length[844]       =   64'h0000000000000100;
assign   tb_i_aad[844]                        =   tb_i_aad[843];
assign   tb_i_rf_static_plaintext_length[844] =   64'h0000000000000280;
assign   tb_i_plaintext[844]                  =   tb_i_plaintext[843];
assign   tb_o_valid[844]                      =   1'b0;
assign   tb_o_sop[844]                        =   1'b0;
assign   tb_o_ciphertext[844]                 =   tb_o_ciphertext[843];
assign   tb_o_tag_ready[844]                  =   1'b0;
assign   tb_o_tag[844]                        =   tb_o_tag[843];

// CLK no. 845/1240
// *************************************************
assign   tb_i_valid[845]                      =   1'b0;
assign   tb_i_reset[845]                      =   1'b0;
assign   tb_i_sop[845]                        =   1'b0;
assign   tb_i_key_update[845]                 =   1'b0;
assign   tb_i_key[845]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[845]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[845]               =   1'b0;
assign   tb_i_rf_static_encrypt[845]          =   1'b1;
assign   tb_i_clear_fault_flags[845]          =   1'b0;
assign   tb_i_rf_static_aad_length[845]       =   64'h0000000000000100;
assign   tb_i_aad[845]                        =   tb_i_aad[844];
assign   tb_i_rf_static_plaintext_length[845] =   64'h0000000000000280;
assign   tb_i_plaintext[845]                  =   tb_i_plaintext[844];
assign   tb_o_valid[845]                      =   1'b0;
assign   tb_o_sop[845]                        =   1'b0;
assign   tb_o_ciphertext[845]                 =   tb_o_ciphertext[844];
assign   tb_o_tag_ready[845]                  =   1'b0;
assign   tb_o_tag[845]                        =   tb_o_tag[844];

// CLK no. 846/1240
// *************************************************
assign   tb_i_valid[846]                      =   1'b0;
assign   tb_i_reset[846]                      =   1'b0;
assign   tb_i_sop[846]                        =   1'b0;
assign   tb_i_key_update[846]                 =   1'b0;
assign   tb_i_key[846]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[846]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[846]               =   1'b0;
assign   tb_i_rf_static_encrypt[846]          =   1'b1;
assign   tb_i_clear_fault_flags[846]          =   1'b0;
assign   tb_i_rf_static_aad_length[846]       =   64'h0000000000000100;
assign   tb_i_aad[846]                        =   tb_i_aad[845];
assign   tb_i_rf_static_plaintext_length[846] =   64'h0000000000000280;
assign   tb_i_plaintext[846]                  =   tb_i_plaintext[845];
assign   tb_o_valid[846]                      =   1'b0;
assign   tb_o_sop[846]                        =   1'b0;
assign   tb_o_ciphertext[846]                 =   tb_o_ciphertext[845];
assign   tb_o_tag_ready[846]                  =   1'b0;
assign   tb_o_tag[846]                        =   tb_o_tag[845];

// CLK no. 847/1240
// *************************************************
assign   tb_i_valid[847]                      =   1'b0;
assign   tb_i_reset[847]                      =   1'b0;
assign   tb_i_sop[847]                        =   1'b0;
assign   tb_i_key_update[847]                 =   1'b0;
assign   tb_i_key[847]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[847]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[847]               =   1'b0;
assign   tb_i_rf_static_encrypt[847]          =   1'b1;
assign   tb_i_clear_fault_flags[847]          =   1'b0;
assign   tb_i_rf_static_aad_length[847]       =   64'h0000000000000100;
assign   tb_i_aad[847]                        =   tb_i_aad[846];
assign   tb_i_rf_static_plaintext_length[847] =   64'h0000000000000280;
assign   tb_i_plaintext[847]                  =   tb_i_plaintext[846];
assign   tb_o_valid[847]                      =   1'b0;
assign   tb_o_sop[847]                        =   1'b0;
assign   tb_o_ciphertext[847]                 =   tb_o_ciphertext[846];
assign   tb_o_tag_ready[847]                  =   1'b0;
assign   tb_o_tag[847]                        =   tb_o_tag[846];

// CLK no. 848/1240
// *************************************************
assign   tb_i_valid[848]                      =   1'b0;
assign   tb_i_reset[848]                      =   1'b0;
assign   tb_i_sop[848]                        =   1'b0;
assign   tb_i_key_update[848]                 =   1'b0;
assign   tb_i_key[848]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[848]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[848]               =   1'b0;
assign   tb_i_rf_static_encrypt[848]          =   1'b1;
assign   tb_i_clear_fault_flags[848]          =   1'b0;
assign   tb_i_rf_static_aad_length[848]       =   64'h0000000000000100;
assign   tb_i_aad[848]                        =   tb_i_aad[847];
assign   tb_i_rf_static_plaintext_length[848] =   64'h0000000000000280;
assign   tb_i_plaintext[848]                  =   tb_i_plaintext[847];
assign   tb_o_valid[848]                      =   1'b0;
assign   tb_o_sop[848]                        =   1'b0;
assign   tb_o_ciphertext[848]                 =   tb_o_ciphertext[847];
assign   tb_o_tag_ready[848]                  =   1'b0;
assign   tb_o_tag[848]                        =   tb_o_tag[847];

// CLK no. 849/1240
// *************************************************
assign   tb_i_valid[849]                      =   1'b0;
assign   tb_i_reset[849]                      =   1'b0;
assign   tb_i_sop[849]                        =   1'b0;
assign   tb_i_key_update[849]                 =   1'b0;
assign   tb_i_key[849]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[849]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[849]               =   1'b0;
assign   tb_i_rf_static_encrypt[849]          =   1'b1;
assign   tb_i_clear_fault_flags[849]          =   1'b0;
assign   tb_i_rf_static_aad_length[849]       =   64'h0000000000000100;
assign   tb_i_aad[849]                        =   tb_i_aad[848];
assign   tb_i_rf_static_plaintext_length[849] =   64'h0000000000000280;
assign   tb_i_plaintext[849]                  =   tb_i_plaintext[848];
assign   tb_o_valid[849]                      =   1'b0;
assign   tb_o_sop[849]                        =   1'b0;
assign   tb_o_ciphertext[849]                 =   tb_o_ciphertext[848];
assign   tb_o_tag_ready[849]                  =   1'b0;
assign   tb_o_tag[849]                        =   tb_o_tag[848];

// CLK no. 850/1240
// *************************************************
assign   tb_i_valid[850]                      =   1'b0;
assign   tb_i_reset[850]                      =   1'b0;
assign   tb_i_sop[850]                        =   1'b0;
assign   tb_i_key_update[850]                 =   1'b0;
assign   tb_i_key[850]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[850]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[850]               =   1'b0;
assign   tb_i_rf_static_encrypt[850]          =   1'b1;
assign   tb_i_clear_fault_flags[850]          =   1'b0;
assign   tb_i_rf_static_aad_length[850]       =   64'h0000000000000100;
assign   tb_i_aad[850]                        =   tb_i_aad[849];
assign   tb_i_rf_static_plaintext_length[850] =   64'h0000000000000280;
assign   tb_i_plaintext[850]                  =   tb_i_plaintext[849];
assign   tb_o_valid[850]                      =   1'b0;
assign   tb_o_sop[850]                        =   1'b0;
assign   tb_o_ciphertext[850]                 =   tb_o_ciphertext[849];
assign   tb_o_tag_ready[850]                  =   1'b0;
assign   tb_o_tag[850]                        =   tb_o_tag[849];

// CLK no. 851/1240
// *************************************************
assign   tb_i_valid[851]                      =   1'b0;
assign   tb_i_reset[851]                      =   1'b0;
assign   tb_i_sop[851]                        =   1'b0;
assign   tb_i_key_update[851]                 =   1'b0;
assign   tb_i_key[851]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[851]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[851]               =   1'b0;
assign   tb_i_rf_static_encrypt[851]          =   1'b1;
assign   tb_i_clear_fault_flags[851]          =   1'b0;
assign   tb_i_rf_static_aad_length[851]       =   64'h0000000000000100;
assign   tb_i_aad[851]                        =   tb_i_aad[850];
assign   tb_i_rf_static_plaintext_length[851] =   64'h0000000000000280;
assign   tb_i_plaintext[851]                  =   tb_i_plaintext[850];
assign   tb_o_valid[851]                      =   1'b0;
assign   tb_o_sop[851]                        =   1'b0;
assign   tb_o_ciphertext[851]                 =   tb_o_ciphertext[850];
assign   tb_o_tag_ready[851]                  =   1'b0;
assign   tb_o_tag[851]                        =   tb_o_tag[850];

// CLK no. 852/1240
// *************************************************
assign   tb_i_valid[852]                      =   1'b0;
assign   tb_i_reset[852]                      =   1'b0;
assign   tb_i_sop[852]                        =   1'b0;
assign   tb_i_key_update[852]                 =   1'b0;
assign   tb_i_key[852]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[852]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[852]               =   1'b0;
assign   tb_i_rf_static_encrypt[852]          =   1'b1;
assign   tb_i_clear_fault_flags[852]          =   1'b0;
assign   tb_i_rf_static_aad_length[852]       =   64'h0000000000000100;
assign   tb_i_aad[852]                        =   tb_i_aad[851];
assign   tb_i_rf_static_plaintext_length[852] =   64'h0000000000000280;
assign   tb_i_plaintext[852]                  =   tb_i_plaintext[851];
assign   tb_o_valid[852]                      =   1'b0;
assign   tb_o_sop[852]                        =   1'b0;
assign   tb_o_ciphertext[852]                 =   tb_o_ciphertext[851];
assign   tb_o_tag_ready[852]                  =   1'b0;
assign   tb_o_tag[852]                        =   tb_o_tag[851];

// CLK no. 853/1240
// *************************************************
assign   tb_i_valid[853]                      =   1'b0;
assign   tb_i_reset[853]                      =   1'b0;
assign   tb_i_sop[853]                        =   1'b0;
assign   tb_i_key_update[853]                 =   1'b0;
assign   tb_i_key[853]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[853]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[853]               =   1'b0;
assign   tb_i_rf_static_encrypt[853]          =   1'b1;
assign   tb_i_clear_fault_flags[853]          =   1'b0;
assign   tb_i_rf_static_aad_length[853]       =   64'h0000000000000100;
assign   tb_i_aad[853]                        =   tb_i_aad[852];
assign   tb_i_rf_static_plaintext_length[853] =   64'h0000000000000280;
assign   tb_i_plaintext[853]                  =   tb_i_plaintext[852];
assign   tb_o_valid[853]                      =   1'b0;
assign   tb_o_sop[853]                        =   1'b0;
assign   tb_o_ciphertext[853]                 =   tb_o_ciphertext[852];
assign   tb_o_tag_ready[853]                  =   1'b0;
assign   tb_o_tag[853]                        =   tb_o_tag[852];

// CLK no. 854/1240
// *************************************************
assign   tb_i_valid[854]                      =   1'b0;
assign   tb_i_reset[854]                      =   1'b0;
assign   tb_i_sop[854]                        =   1'b0;
assign   tb_i_key_update[854]                 =   1'b0;
assign   tb_i_key[854]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[854]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[854]               =   1'b0;
assign   tb_i_rf_static_encrypt[854]          =   1'b1;
assign   tb_i_clear_fault_flags[854]          =   1'b0;
assign   tb_i_rf_static_aad_length[854]       =   64'h0000000000000100;
assign   tb_i_aad[854]                        =   tb_i_aad[853];
assign   tb_i_rf_static_plaintext_length[854] =   64'h0000000000000280;
assign   tb_i_plaintext[854]                  =   tb_i_plaintext[853];
assign   tb_o_valid[854]                      =   1'b0;
assign   tb_o_sop[854]                        =   1'b0;
assign   tb_o_ciphertext[854]                 =   tb_o_ciphertext[853];
assign   tb_o_tag_ready[854]                  =   1'b0;
assign   tb_o_tag[854]                        =   tb_o_tag[853];

// CLK no. 855/1240
// *************************************************
assign   tb_i_valid[855]                      =   1'b0;
assign   tb_i_reset[855]                      =   1'b0;
assign   tb_i_sop[855]                        =   1'b0;
assign   tb_i_key_update[855]                 =   1'b0;
assign   tb_i_key[855]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[855]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[855]               =   1'b0;
assign   tb_i_rf_static_encrypt[855]          =   1'b1;
assign   tb_i_clear_fault_flags[855]          =   1'b0;
assign   tb_i_rf_static_aad_length[855]       =   64'h0000000000000100;
assign   tb_i_aad[855]                        =   tb_i_aad[854];
assign   tb_i_rf_static_plaintext_length[855] =   64'h0000000000000280;
assign   tb_i_plaintext[855]                  =   tb_i_plaintext[854];
assign   tb_o_valid[855]                      =   1'b0;
assign   tb_o_sop[855]                        =   1'b0;
assign   tb_o_ciphertext[855]                 =   tb_o_ciphertext[854];
assign   tb_o_tag_ready[855]                  =   1'b0;
assign   tb_o_tag[855]                        =   tb_o_tag[854];

// CLK no. 856/1240
// *************************************************
assign   tb_i_valid[856]                      =   1'b0;
assign   tb_i_reset[856]                      =   1'b0;
assign   tb_i_sop[856]                        =   1'b0;
assign   tb_i_key_update[856]                 =   1'b0;
assign   tb_i_key[856]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[856]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[856]               =   1'b0;
assign   tb_i_rf_static_encrypt[856]          =   1'b1;
assign   tb_i_clear_fault_flags[856]          =   1'b0;
assign   tb_i_rf_static_aad_length[856]       =   64'h0000000000000100;
assign   tb_i_aad[856]                        =   tb_i_aad[855];
assign   tb_i_rf_static_plaintext_length[856] =   64'h0000000000000280;
assign   tb_i_plaintext[856]                  =   tb_i_plaintext[855];
assign   tb_o_valid[856]                      =   1'b0;
assign   tb_o_sop[856]                        =   1'b0;
assign   tb_o_ciphertext[856]                 =   tb_o_ciphertext[855];
assign   tb_o_tag_ready[856]                  =   1'b0;
assign   tb_o_tag[856]                        =   tb_o_tag[855];

// CLK no. 857/1240
// *************************************************
assign   tb_i_valid[857]                      =   1'b0;
assign   tb_i_reset[857]                      =   1'b0;
assign   tb_i_sop[857]                        =   1'b0;
assign   tb_i_key_update[857]                 =   1'b0;
assign   tb_i_key[857]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[857]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[857]               =   1'b0;
assign   tb_i_rf_static_encrypt[857]          =   1'b1;
assign   tb_i_clear_fault_flags[857]          =   1'b0;
assign   tb_i_rf_static_aad_length[857]       =   64'h0000000000000100;
assign   tb_i_aad[857]                        =   tb_i_aad[856];
assign   tb_i_rf_static_plaintext_length[857] =   64'h0000000000000280;
assign   tb_i_plaintext[857]                  =   tb_i_plaintext[856];
assign   tb_o_valid[857]                      =   1'b0;
assign   tb_o_sop[857]                        =   1'b0;
assign   tb_o_ciphertext[857]                 =   tb_o_ciphertext[856];
assign   tb_o_tag_ready[857]                  =   1'b0;
assign   tb_o_tag[857]                        =   tb_o_tag[856];

// CLK no. 858/1240
// *************************************************
assign   tb_i_valid[858]                      =   1'b0;
assign   tb_i_reset[858]                      =   1'b0;
assign   tb_i_sop[858]                        =   1'b0;
assign   tb_i_key_update[858]                 =   1'b0;
assign   tb_i_key[858]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[858]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[858]               =   1'b0;
assign   tb_i_rf_static_encrypt[858]          =   1'b1;
assign   tb_i_clear_fault_flags[858]          =   1'b0;
assign   tb_i_rf_static_aad_length[858]       =   64'h0000000000000100;
assign   tb_i_aad[858]                        =   tb_i_aad[857];
assign   tb_i_rf_static_plaintext_length[858] =   64'h0000000000000280;
assign   tb_i_plaintext[858]                  =   tb_i_plaintext[857];
assign   tb_o_valid[858]                      =   1'b0;
assign   tb_o_sop[858]                        =   1'b0;
assign   tb_o_ciphertext[858]                 =   tb_o_ciphertext[857];
assign   tb_o_tag_ready[858]                  =   1'b0;
assign   tb_o_tag[858]                        =   tb_o_tag[857];

// CLK no. 859/1240
// *************************************************
assign   tb_i_valid[859]                      =   1'b0;
assign   tb_i_reset[859]                      =   1'b0;
assign   tb_i_sop[859]                        =   1'b0;
assign   tb_i_key_update[859]                 =   1'b0;
assign   tb_i_key[859]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[859]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[859]               =   1'b0;
assign   tb_i_rf_static_encrypt[859]          =   1'b1;
assign   tb_i_clear_fault_flags[859]          =   1'b0;
assign   tb_i_rf_static_aad_length[859]       =   64'h0000000000000100;
assign   tb_i_aad[859]                        =   tb_i_aad[858];
assign   tb_i_rf_static_plaintext_length[859] =   64'h0000000000000280;
assign   tb_i_plaintext[859]                  =   tb_i_plaintext[858];
assign   tb_o_valid[859]                      =   1'b0;
assign   tb_o_sop[859]                        =   1'b0;
assign   tb_o_ciphertext[859]                 =   tb_o_ciphertext[858];
assign   tb_o_tag_ready[859]                  =   1'b0;
assign   tb_o_tag[859]                        =   tb_o_tag[858];

// CLK no. 860/1240
// *************************************************
assign   tb_i_valid[860]                      =   1'b0;
assign   tb_i_reset[860]                      =   1'b0;
assign   tb_i_sop[860]                        =   1'b0;
assign   tb_i_key_update[860]                 =   1'b0;
assign   tb_i_key[860]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[860]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[860]               =   1'b0;
assign   tb_i_rf_static_encrypt[860]          =   1'b1;
assign   tb_i_clear_fault_flags[860]          =   1'b0;
assign   tb_i_rf_static_aad_length[860]       =   64'h0000000000000100;
assign   tb_i_aad[860]                        =   tb_i_aad[859];
assign   tb_i_rf_static_plaintext_length[860] =   64'h0000000000000280;
assign   tb_i_plaintext[860]                  =   tb_i_plaintext[859];
assign   tb_o_valid[860]                      =   1'b0;
assign   tb_o_sop[860]                        =   1'b0;
assign   tb_o_ciphertext[860]                 =   tb_o_ciphertext[859];
assign   tb_o_tag_ready[860]                  =   1'b0;
assign   tb_o_tag[860]                        =   tb_o_tag[859];

// CLK no. 861/1240
// *************************************************
assign   tb_i_valid[861]                      =   1'b0;
assign   tb_i_reset[861]                      =   1'b0;
assign   tb_i_sop[861]                        =   1'b0;
assign   tb_i_key_update[861]                 =   1'b0;
assign   tb_i_key[861]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[861]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[861]               =   1'b0;
assign   tb_i_rf_static_encrypt[861]          =   1'b1;
assign   tb_i_clear_fault_flags[861]          =   1'b0;
assign   tb_i_rf_static_aad_length[861]       =   64'h0000000000000100;
assign   tb_i_aad[861]                        =   tb_i_aad[860];
assign   tb_i_rf_static_plaintext_length[861] =   64'h0000000000000280;
assign   tb_i_plaintext[861]                  =   tb_i_plaintext[860];
assign   tb_o_valid[861]                      =   1'b0;
assign   tb_o_sop[861]                        =   1'b0;
assign   tb_o_ciphertext[861]                 =   tb_o_ciphertext[860];
assign   tb_o_tag_ready[861]                  =   1'b0;
assign   tb_o_tag[861]                        =   tb_o_tag[860];

// CLK no. 862/1240
// *************************************************
assign   tb_i_valid[862]                      =   1'b0;
assign   tb_i_reset[862]                      =   1'b0;
assign   tb_i_sop[862]                        =   1'b0;
assign   tb_i_key_update[862]                 =   1'b0;
assign   tb_i_key[862]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[862]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[862]               =   1'b0;
assign   tb_i_rf_static_encrypt[862]          =   1'b1;
assign   tb_i_clear_fault_flags[862]          =   1'b0;
assign   tb_i_rf_static_aad_length[862]       =   64'h0000000000000100;
assign   tb_i_aad[862]                        =   tb_i_aad[861];
assign   tb_i_rf_static_plaintext_length[862] =   64'h0000000000000280;
assign   tb_i_plaintext[862]                  =   tb_i_plaintext[861];
assign   tb_o_valid[862]                      =   1'b0;
assign   tb_o_sop[862]                        =   1'b0;
assign   tb_o_ciphertext[862]                 =   tb_o_ciphertext[861];
assign   tb_o_tag_ready[862]                  =   1'b0;
assign   tb_o_tag[862]                        =   tb_o_tag[861];

// CLK no. 863/1240
// *************************************************
assign   tb_i_valid[863]                      =   1'b0;
assign   tb_i_reset[863]                      =   1'b0;
assign   tb_i_sop[863]                        =   1'b0;
assign   tb_i_key_update[863]                 =   1'b0;
assign   tb_i_key[863]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[863]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[863]               =   1'b0;
assign   tb_i_rf_static_encrypt[863]          =   1'b1;
assign   tb_i_clear_fault_flags[863]          =   1'b0;
assign   tb_i_rf_static_aad_length[863]       =   64'h0000000000000100;
assign   tb_i_aad[863]                        =   tb_i_aad[862];
assign   tb_i_rf_static_plaintext_length[863] =   64'h0000000000000280;
assign   tb_i_plaintext[863]                  =   tb_i_plaintext[862];
assign   tb_o_valid[863]                      =   1'b0;
assign   tb_o_sop[863]                        =   1'b0;
assign   tb_o_ciphertext[863]                 =   tb_o_ciphertext[862];
assign   tb_o_tag_ready[863]                  =   1'b0;
assign   tb_o_tag[863]                        =   tb_o_tag[862];

// CLK no. 864/1240
// *************************************************
assign   tb_i_valid[864]                      =   1'b0;
assign   tb_i_reset[864]                      =   1'b0;
assign   tb_i_sop[864]                        =   1'b0;
assign   tb_i_key_update[864]                 =   1'b0;
assign   tb_i_key[864]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[864]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[864]               =   1'b0;
assign   tb_i_rf_static_encrypt[864]          =   1'b1;
assign   tb_i_clear_fault_flags[864]          =   1'b0;
assign   tb_i_rf_static_aad_length[864]       =   64'h0000000000000100;
assign   tb_i_aad[864]                        =   tb_i_aad[863];
assign   tb_i_rf_static_plaintext_length[864] =   64'h0000000000000280;
assign   tb_i_plaintext[864]                  =   tb_i_plaintext[863];
assign   tb_o_valid[864]                      =   1'b0;
assign   tb_o_sop[864]                        =   1'b0;
assign   tb_o_ciphertext[864]                 =   tb_o_ciphertext[863];
assign   tb_o_tag_ready[864]                  =   1'b0;
assign   tb_o_tag[864]                        =   tb_o_tag[863];

// CLK no. 865/1240
// *************************************************
assign   tb_i_valid[865]                      =   1'b0;
assign   tb_i_reset[865]                      =   1'b0;
assign   tb_i_sop[865]                        =   1'b0;
assign   tb_i_key_update[865]                 =   1'b0;
assign   tb_i_key[865]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[865]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[865]               =   1'b0;
assign   tb_i_rf_static_encrypt[865]          =   1'b1;
assign   tb_i_clear_fault_flags[865]          =   1'b0;
assign   tb_i_rf_static_aad_length[865]       =   64'h0000000000000100;
assign   tb_i_aad[865]                        =   tb_i_aad[864];
assign   tb_i_rf_static_plaintext_length[865] =   64'h0000000000000280;
assign   tb_i_plaintext[865]                  =   tb_i_plaintext[864];
assign   tb_o_valid[865]                      =   1'b0;
assign   tb_o_sop[865]                        =   1'b0;
assign   tb_o_ciphertext[865]                 =   tb_o_ciphertext[864];
assign   tb_o_tag_ready[865]                  =   1'b0;
assign   tb_o_tag[865]                        =   tb_o_tag[864];

// CLK no. 866/1240
// *************************************************
assign   tb_i_valid[866]                      =   1'b0;
assign   tb_i_reset[866]                      =   1'b0;
assign   tb_i_sop[866]                        =   1'b0;
assign   tb_i_key_update[866]                 =   1'b0;
assign   tb_i_key[866]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[866]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[866]               =   1'b0;
assign   tb_i_rf_static_encrypt[866]          =   1'b1;
assign   tb_i_clear_fault_flags[866]          =   1'b0;
assign   tb_i_rf_static_aad_length[866]       =   64'h0000000000000100;
assign   tb_i_aad[866]                        =   tb_i_aad[865];
assign   tb_i_rf_static_plaintext_length[866] =   64'h0000000000000280;
assign   tb_i_plaintext[866]                  =   tb_i_plaintext[865];
assign   tb_o_valid[866]                      =   1'b0;
assign   tb_o_sop[866]                        =   1'b0;
assign   tb_o_ciphertext[866]                 =   tb_o_ciphertext[865];
assign   tb_o_tag_ready[866]                  =   1'b0;
assign   tb_o_tag[866]                        =   tb_o_tag[865];

// CLK no. 867/1240
// *************************************************
assign   tb_i_valid[867]                      =   1'b0;
assign   tb_i_reset[867]                      =   1'b0;
assign   tb_i_sop[867]                        =   1'b0;
assign   tb_i_key_update[867]                 =   1'b0;
assign   tb_i_key[867]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[867]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[867]               =   1'b0;
assign   tb_i_rf_static_encrypt[867]          =   1'b1;
assign   tb_i_clear_fault_flags[867]          =   1'b0;
assign   tb_i_rf_static_aad_length[867]       =   64'h0000000000000100;
assign   tb_i_aad[867]                        =   tb_i_aad[866];
assign   tb_i_rf_static_plaintext_length[867] =   64'h0000000000000280;
assign   tb_i_plaintext[867]                  =   tb_i_plaintext[866];
assign   tb_o_valid[867]                      =   1'b0;
assign   tb_o_sop[867]                        =   1'b0;
assign   tb_o_ciphertext[867]                 =   tb_o_ciphertext[866];
assign   tb_o_tag_ready[867]                  =   1'b0;
assign   tb_o_tag[867]                        =   tb_o_tag[866];

// CLK no. 868/1240
// *************************************************
assign   tb_i_valid[868]                      =   1'b0;
assign   tb_i_reset[868]                      =   1'b0;
assign   tb_i_sop[868]                        =   1'b0;
assign   tb_i_key_update[868]                 =   1'b0;
assign   tb_i_key[868]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[868]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[868]               =   1'b0;
assign   tb_i_rf_static_encrypt[868]          =   1'b1;
assign   tb_i_clear_fault_flags[868]          =   1'b0;
assign   tb_i_rf_static_aad_length[868]       =   64'h0000000000000100;
assign   tb_i_aad[868]                        =   tb_i_aad[867];
assign   tb_i_rf_static_plaintext_length[868] =   64'h0000000000000280;
assign   tb_i_plaintext[868]                  =   tb_i_plaintext[867];
assign   tb_o_valid[868]                      =   1'b0;
assign   tb_o_sop[868]                        =   1'b0;
assign   tb_o_ciphertext[868]                 =   tb_o_ciphertext[867];
assign   tb_o_tag_ready[868]                  =   1'b0;
assign   tb_o_tag[868]                        =   tb_o_tag[867];

// CLK no. 869/1240
// *************************************************
assign   tb_i_valid[869]                      =   1'b0;
assign   tb_i_reset[869]                      =   1'b0;
assign   tb_i_sop[869]                        =   1'b0;
assign   tb_i_key_update[869]                 =   1'b0;
assign   tb_i_key[869]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[869]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[869]               =   1'b0;
assign   tb_i_rf_static_encrypt[869]          =   1'b1;
assign   tb_i_clear_fault_flags[869]          =   1'b0;
assign   tb_i_rf_static_aad_length[869]       =   64'h0000000000000100;
assign   tb_i_aad[869]                        =   tb_i_aad[868];
assign   tb_i_rf_static_plaintext_length[869] =   64'h0000000000000280;
assign   tb_i_plaintext[869]                  =   tb_i_plaintext[868];
assign   tb_o_valid[869]                      =   1'b0;
assign   tb_o_sop[869]                        =   1'b0;
assign   tb_o_ciphertext[869]                 =   tb_o_ciphertext[868];
assign   tb_o_tag_ready[869]                  =   1'b0;
assign   tb_o_tag[869]                        =   tb_o_tag[868];

// CLK no. 870/1240
// *************************************************
assign   tb_i_valid[870]                      =   1'b0;
assign   tb_i_reset[870]                      =   1'b0;
assign   tb_i_sop[870]                        =   1'b0;
assign   tb_i_key_update[870]                 =   1'b0;
assign   tb_i_key[870]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[870]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[870]               =   1'b0;
assign   tb_i_rf_static_encrypt[870]          =   1'b1;
assign   tb_i_clear_fault_flags[870]          =   1'b0;
assign   tb_i_rf_static_aad_length[870]       =   64'h0000000000000100;
assign   tb_i_aad[870]                        =   tb_i_aad[869];
assign   tb_i_rf_static_plaintext_length[870] =   64'h0000000000000280;
assign   tb_i_plaintext[870]                  =   tb_i_plaintext[869];
assign   tb_o_valid[870]                      =   1'b0;
assign   tb_o_sop[870]                        =   1'b0;
assign   tb_o_ciphertext[870]                 =   tb_o_ciphertext[869];
assign   tb_o_tag_ready[870]                  =   1'b0;
assign   tb_o_tag[870]                        =   tb_o_tag[869];

// CLK no. 871/1240
// *************************************************
assign   tb_i_valid[871]                      =   1'b0;
assign   tb_i_reset[871]                      =   1'b0;
assign   tb_i_sop[871]                        =   1'b0;
assign   tb_i_key_update[871]                 =   1'b0;
assign   tb_i_key[871]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[871]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[871]               =   1'b0;
assign   tb_i_rf_static_encrypt[871]          =   1'b1;
assign   tb_i_clear_fault_flags[871]          =   1'b0;
assign   tb_i_rf_static_aad_length[871]       =   64'h0000000000000100;
assign   tb_i_aad[871]                        =   tb_i_aad[870];
assign   tb_i_rf_static_plaintext_length[871] =   64'h0000000000000280;
assign   tb_i_plaintext[871]                  =   tb_i_plaintext[870];
assign   tb_o_valid[871]                      =   1'b0;
assign   tb_o_sop[871]                        =   1'b0;
assign   tb_o_ciphertext[871]                 =   tb_o_ciphertext[870];
assign   tb_o_tag_ready[871]                  =   1'b0;
assign   tb_o_tag[871]                        =   tb_o_tag[870];

// CLK no. 872/1240
// *************************************************
assign   tb_i_valid[872]                      =   1'b0;
assign   tb_i_reset[872]                      =   1'b0;
assign   tb_i_sop[872]                        =   1'b0;
assign   tb_i_key_update[872]                 =   1'b0;
assign   tb_i_key[872]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[872]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[872]               =   1'b0;
assign   tb_i_rf_static_encrypt[872]          =   1'b1;
assign   tb_i_clear_fault_flags[872]          =   1'b0;
assign   tb_i_rf_static_aad_length[872]       =   64'h0000000000000100;
assign   tb_i_aad[872]                        =   tb_i_aad[871];
assign   tb_i_rf_static_plaintext_length[872] =   64'h0000000000000280;
assign   tb_i_plaintext[872]                  =   tb_i_plaintext[871];
assign   tb_o_valid[872]                      =   1'b0;
assign   tb_o_sop[872]                        =   1'b0;
assign   tb_o_ciphertext[872]                 =   tb_o_ciphertext[871];
assign   tb_o_tag_ready[872]                  =   1'b0;
assign   tb_o_tag[872]                        =   tb_o_tag[871];

// CLK no. 873/1240
// *************************************************
assign   tb_i_valid[873]                      =   1'b0;
assign   tb_i_reset[873]                      =   1'b0;
assign   tb_i_sop[873]                        =   1'b0;
assign   tb_i_key_update[873]                 =   1'b0;
assign   tb_i_key[873]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[873]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[873]               =   1'b0;
assign   tb_i_rf_static_encrypt[873]          =   1'b1;
assign   tb_i_clear_fault_flags[873]          =   1'b0;
assign   tb_i_rf_static_aad_length[873]       =   64'h0000000000000100;
assign   tb_i_aad[873]                        =   tb_i_aad[872];
assign   tb_i_rf_static_plaintext_length[873] =   64'h0000000000000280;
assign   tb_i_plaintext[873]                  =   tb_i_plaintext[872];
assign   tb_o_valid[873]                      =   1'b1;
assign   tb_o_sop[873]                        =   1'b1;
assign   tb_o_ciphertext[873]                 =   256'h9be2b568a654952541a82a15e0cef5c8a43dacbef6efb4e596eba46733555c0f;
assign   tb_o_tag_ready[873]                  =   1'b0;
assign   tb_o_tag[873]                        =   tb_o_tag[872];

// CLK no. 874/1240
// *************************************************
assign   tb_i_valid[874]                      =   1'b0;
assign   tb_i_reset[874]                      =   1'b0;
assign   tb_i_sop[874]                        =   1'b0;
assign   tb_i_key_update[874]                 =   1'b0;
assign   tb_i_key[874]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[874]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[874]               =   1'b0;
assign   tb_i_rf_static_encrypt[874]          =   1'b1;
assign   tb_i_clear_fault_flags[874]          =   1'b0;
assign   tb_i_rf_static_aad_length[874]       =   64'h0000000000000100;
assign   tb_i_aad[874]                        =   tb_i_aad[873];
assign   tb_i_rf_static_plaintext_length[874] =   64'h0000000000000280;
assign   tb_i_plaintext[874]                  =   tb_i_plaintext[873];
assign   tb_o_valid[874]                      =   1'b1;
assign   tb_o_sop[874]                        =   1'b0;
assign   tb_o_ciphertext[874]                 =   256'hfdd3e685726155d1f7ec8c58d4b566c4cbef31b80486aa4b8e54eb4adfdabfc6;
assign   tb_o_tag_ready[874]                  =   1'b0;
assign   tb_o_tag[874]                        =   tb_o_tag[873];

// CLK no. 875/1240
// *************************************************
assign   tb_i_valid[875]                      =   1'b0;
assign   tb_i_reset[875]                      =   1'b0;
assign   tb_i_sop[875]                        =   1'b0;
assign   tb_i_key_update[875]                 =   1'b0;
assign   tb_i_key[875]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[875]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[875]               =   1'b0;
assign   tb_i_rf_static_encrypt[875]          =   1'b1;
assign   tb_i_clear_fault_flags[875]          =   1'b0;
assign   tb_i_rf_static_aad_length[875]       =   64'h0000000000000100;
assign   tb_i_aad[875]                        =   tb_i_aad[874];
assign   tb_i_rf_static_plaintext_length[875] =   64'h0000000000000280;
assign   tb_i_plaintext[875]                  =   tb_i_plaintext[874];
assign   tb_o_valid[875]                      =   1'b1;
assign   tb_o_sop[875]                        =   1'b0;
assign   tb_o_ciphertext[875]                 =   256'he028fe2b7b0a0b0ce2281f34d714e5fc;
assign   tb_o_tag_ready[875]                  =   1'b0;
assign   tb_o_tag[875]                        =   tb_o_tag[874];

// CLK no. 876/1240
// *************************************************
assign   tb_i_valid[876]                      =   1'b0;
assign   tb_i_reset[876]                      =   1'b0;
assign   tb_i_sop[876]                        =   1'b0;
assign   tb_i_key_update[876]                 =   1'b0;
assign   tb_i_key[876]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[876]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[876]               =   1'b0;
assign   tb_i_rf_static_encrypt[876]          =   1'b1;
assign   tb_i_clear_fault_flags[876]          =   1'b0;
assign   tb_i_rf_static_aad_length[876]       =   64'h0000000000000100;
assign   tb_i_aad[876]                        =   tb_i_aad[875];
assign   tb_i_rf_static_plaintext_length[876] =   64'h0000000000000280;
assign   tb_i_plaintext[876]                  =   tb_i_plaintext[875];
assign   tb_o_valid[876]                      =   1'b0;
assign   tb_o_sop[876]                        =   1'b0;
assign   tb_o_ciphertext[876]                 =   tb_o_ciphertext[875];
assign   tb_o_tag_ready[876]                  =   1'b0;
assign   tb_o_tag[876]                        =   tb_o_tag[875];

// CLK no. 877/1240
// *************************************************
assign   tb_i_valid[877]                      =   1'b0;
assign   tb_i_reset[877]                      =   1'b0;
assign   tb_i_sop[877]                        =   1'b0;
assign   tb_i_key_update[877]                 =   1'b0;
assign   tb_i_key[877]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[877]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[877]               =   1'b0;
assign   tb_i_rf_static_encrypt[877]          =   1'b1;
assign   tb_i_clear_fault_flags[877]          =   1'b0;
assign   tb_i_rf_static_aad_length[877]       =   64'h0000000000000100;
assign   tb_i_aad[877]                        =   tb_i_aad[876];
assign   tb_i_rf_static_plaintext_length[877] =   64'h0000000000000280;
assign   tb_i_plaintext[877]                  =   tb_i_plaintext[876];
assign   tb_o_valid[877]                      =   1'b0;
assign   tb_o_sop[877]                        =   1'b0;
assign   tb_o_ciphertext[877]                 =   tb_o_ciphertext[876];
assign   tb_o_tag_ready[877]                  =   1'b0;
assign   tb_o_tag[877]                        =   tb_o_tag[876];

// CLK no. 878/1240
// *************************************************
assign   tb_i_valid[878]                      =   1'b0;
assign   tb_i_reset[878]                      =   1'b0;
assign   tb_i_sop[878]                        =   1'b0;
assign   tb_i_key_update[878]                 =   1'b0;
assign   tb_i_key[878]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[878]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[878]               =   1'b0;
assign   tb_i_rf_static_encrypt[878]          =   1'b1;
assign   tb_i_clear_fault_flags[878]          =   1'b0;
assign   tb_i_rf_static_aad_length[878]       =   64'h0000000000000100;
assign   tb_i_aad[878]                        =   tb_i_aad[877];
assign   tb_i_rf_static_plaintext_length[878] =   64'h0000000000000280;
assign   tb_i_plaintext[878]                  =   tb_i_plaintext[877];
assign   tb_o_valid[878]                      =   1'b0;
assign   tb_o_sop[878]                        =   1'b0;
assign   tb_o_ciphertext[878]                 =   tb_o_ciphertext[877];
assign   tb_o_tag_ready[878]                  =   1'b0;
assign   tb_o_tag[878]                        =   tb_o_tag[877];

// CLK no. 879/1240
// *************************************************
assign   tb_i_valid[879]                      =   1'b0;
assign   tb_i_reset[879]                      =   1'b0;
assign   tb_i_sop[879]                        =   1'b0;
assign   tb_i_key_update[879]                 =   1'b0;
assign   tb_i_key[879]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[879]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[879]               =   1'b0;
assign   tb_i_rf_static_encrypt[879]          =   1'b1;
assign   tb_i_clear_fault_flags[879]          =   1'b0;
assign   tb_i_rf_static_aad_length[879]       =   64'h0000000000000100;
assign   tb_i_aad[879]                        =   tb_i_aad[878];
assign   tb_i_rf_static_plaintext_length[879] =   64'h0000000000000280;
assign   tb_i_plaintext[879]                  =   tb_i_plaintext[878];
assign   tb_o_valid[879]                      =   1'b0;
assign   tb_o_sop[879]                        =   1'b0;
assign   tb_o_ciphertext[879]                 =   tb_o_ciphertext[878];
assign   tb_o_tag_ready[879]                  =   1'b0;
assign   tb_o_tag[879]                        =   tb_o_tag[878];

// CLK no. 880/1240
// *************************************************
assign   tb_i_valid[880]                      =   1'b0;
assign   tb_i_reset[880]                      =   1'b0;
assign   tb_i_sop[880]                        =   1'b0;
assign   tb_i_key_update[880]                 =   1'b0;
assign   tb_i_key[880]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[880]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[880]               =   1'b0;
assign   tb_i_rf_static_encrypt[880]          =   1'b1;
assign   tb_i_clear_fault_flags[880]          =   1'b0;
assign   tb_i_rf_static_aad_length[880]       =   64'h0000000000000100;
assign   tb_i_aad[880]                        =   tb_i_aad[879];
assign   tb_i_rf_static_plaintext_length[880] =   64'h0000000000000280;
assign   tb_i_plaintext[880]                  =   tb_i_plaintext[879];
assign   tb_o_valid[880]                      =   1'b0;
assign   tb_o_sop[880]                        =   1'b0;
assign   tb_o_ciphertext[880]                 =   tb_o_ciphertext[879];
assign   tb_o_tag_ready[880]                  =   1'b0;
assign   tb_o_tag[880]                        =   tb_o_tag[879];

// CLK no. 881/1240
// *************************************************
assign   tb_i_valid[881]                      =   1'b0;
assign   tb_i_reset[881]                      =   1'b0;
assign   tb_i_sop[881]                        =   1'b0;
assign   tb_i_key_update[881]                 =   1'b0;
assign   tb_i_key[881]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[881]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[881]               =   1'b0;
assign   tb_i_rf_static_encrypt[881]          =   1'b1;
assign   tb_i_clear_fault_flags[881]          =   1'b0;
assign   tb_i_rf_static_aad_length[881]       =   64'h0000000000000100;
assign   tb_i_aad[881]                        =   tb_i_aad[880];
assign   tb_i_rf_static_plaintext_length[881] =   64'h0000000000000280;
assign   tb_i_plaintext[881]                  =   tb_i_plaintext[880];
assign   tb_o_valid[881]                      =   1'b0;
assign   tb_o_sop[881]                        =   1'b0;
assign   tb_o_ciphertext[881]                 =   tb_o_ciphertext[880];
assign   tb_o_tag_ready[881]                  =   1'b0;
assign   tb_o_tag[881]                        =   tb_o_tag[880];

// CLK no. 882/1240
// *************************************************
assign   tb_i_valid[882]                      =   1'b0;
assign   tb_i_reset[882]                      =   1'b0;
assign   tb_i_sop[882]                        =   1'b0;
assign   tb_i_key_update[882]                 =   1'b0;
assign   tb_i_key[882]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[882]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[882]               =   1'b0;
assign   tb_i_rf_static_encrypt[882]          =   1'b1;
assign   tb_i_clear_fault_flags[882]          =   1'b0;
assign   tb_i_rf_static_aad_length[882]       =   64'h0000000000000100;
assign   tb_i_aad[882]                        =   tb_i_aad[881];
assign   tb_i_rf_static_plaintext_length[882] =   64'h0000000000000280;
assign   tb_i_plaintext[882]                  =   tb_i_plaintext[881];
assign   tb_o_valid[882]                      =   1'b0;
assign   tb_o_sop[882]                        =   1'b0;
assign   tb_o_ciphertext[882]                 =   tb_o_ciphertext[881];
assign   tb_o_tag_ready[882]                  =   1'b0;
assign   tb_o_tag[882]                        =   tb_o_tag[881];

// CLK no. 883/1240
// *************************************************
assign   tb_i_valid[883]                      =   1'b0;
assign   tb_i_reset[883]                      =   1'b0;
assign   tb_i_sop[883]                        =   1'b0;
assign   tb_i_key_update[883]                 =   1'b0;
assign   tb_i_key[883]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[883]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[883]               =   1'b0;
assign   tb_i_rf_static_encrypt[883]          =   1'b1;
assign   tb_i_clear_fault_flags[883]          =   1'b0;
assign   tb_i_rf_static_aad_length[883]       =   64'h0000000000000100;
assign   tb_i_aad[883]                        =   tb_i_aad[882];
assign   tb_i_rf_static_plaintext_length[883] =   64'h0000000000000280;
assign   tb_i_plaintext[883]                  =   tb_i_plaintext[882];
assign   tb_o_valid[883]                      =   1'b0;
assign   tb_o_sop[883]                        =   1'b0;
assign   tb_o_ciphertext[883]                 =   tb_o_ciphertext[882];
assign   tb_o_tag_ready[883]                  =   1'b1;
assign   tb_o_tag[883]                        =   128'h8d8778c6988648b2305e5356cedcc9a1;

// CLK no. 884/1240
// *************************************************
assign   tb_i_valid[884]                      =   1'b0;
assign   tb_i_reset[884]                      =   1'b0;
assign   tb_i_sop[884]                        =   1'b0;
assign   tb_i_key_update[884]                 =   1'b0;
assign   tb_i_key[884]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[884]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[884]               =   1'b0;
assign   tb_i_rf_static_encrypt[884]          =   1'b1;
assign   tb_i_clear_fault_flags[884]          =   1'b0;
assign   tb_i_rf_static_aad_length[884]       =   64'h0000000000000100;
assign   tb_i_aad[884]                        =   tb_i_aad[883];
assign   tb_i_rf_static_plaintext_length[884] =   64'h0000000000000280;
assign   tb_i_plaintext[884]                  =   tb_i_plaintext[883];
assign   tb_o_valid[884]                      =   1'b0;
assign   tb_o_sop[884]                        =   1'b0;
assign   tb_o_ciphertext[884]                 =   tb_o_ciphertext[883];
assign   tb_o_tag_ready[884]                  =   1'b0;
assign   tb_o_tag[884]                        =   tb_o_tag[883];

// CLK no. 885/1240
// *************************************************
assign   tb_i_valid[885]                      =   1'b0;
assign   tb_i_reset[885]                      =   1'b0;
assign   tb_i_sop[885]                        =   1'b0;
assign   tb_i_key_update[885]                 =   1'b0;
assign   tb_i_key[885]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[885]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[885]               =   1'b0;
assign   tb_i_rf_static_encrypt[885]          =   1'b1;
assign   tb_i_clear_fault_flags[885]          =   1'b0;
assign   tb_i_rf_static_aad_length[885]       =   64'h0000000000000100;
assign   tb_i_aad[885]                        =   tb_i_aad[884];
assign   tb_i_rf_static_plaintext_length[885] =   64'h0000000000000280;
assign   tb_i_plaintext[885]                  =   tb_i_plaintext[884];
assign   tb_o_valid[885]                      =   1'b0;
assign   tb_o_sop[885]                        =   1'b0;
assign   tb_o_ciphertext[885]                 =   tb_o_ciphertext[884];
assign   tb_o_tag_ready[885]                  =   1'b0;
assign   tb_o_tag[885]                        =   tb_o_tag[884];

// CLK no. 886/1240
// *************************************************
assign   tb_i_valid[886]                      =   1'b0;
assign   tb_i_reset[886]                      =   1'b0;
assign   tb_i_sop[886]                        =   1'b1;
assign   tb_i_key_update[886]                 =   1'b0;
assign   tb_i_key[886]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[886]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[886]               =   1'b0;
assign   tb_i_rf_static_encrypt[886]          =   1'b1;
assign   tb_i_clear_fault_flags[886]          =   1'b0;
assign   tb_i_rf_static_aad_length[886]       =   64'h0000000000000100;
assign   tb_i_aad[886]                        =   tb_i_aad[885];
assign   tb_i_rf_static_plaintext_length[886] =   64'h0000000000000280;
assign   tb_i_plaintext[886]                  =   tb_i_plaintext[885];
assign   tb_o_valid[886]                      =   1'b0;
assign   tb_o_sop[886]                        =   1'b0;
assign   tb_o_ciphertext[886]                 =   tb_o_ciphertext[885];
assign   tb_o_tag_ready[886]                  =   1'b0;
assign   tb_o_tag[886]                        =   tb_o_tag[885];

// CLK no. 887/1240
// *************************************************
assign   tb_i_valid[887]                      =   1'b1;
assign   tb_i_reset[887]                      =   1'b0;
assign   tb_i_sop[887]                        =   1'b0;
assign   tb_i_key_update[887]                 =   1'b0;
assign   tb_i_key[887]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[887]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[887]               =   1'b0;
assign   tb_i_rf_static_encrypt[887]          =   1'b1;
assign   tb_i_clear_fault_flags[887]          =   1'b0;
assign   tb_i_rf_static_aad_length[887]       =   64'h0000000000000100;
assign   tb_i_aad[887]                        =   256'hc8c1e50584ee8f3948880ba725f7f7b847b584ace67a36f932a4a64228cdf880;
assign   tb_i_rf_static_plaintext_length[887] =   64'h0000000000000280;
assign   tb_i_plaintext[887]                  =   tb_i_plaintext[886];
assign   tb_o_valid[887]                      =   1'b0;
assign   tb_o_sop[887]                        =   1'b0;
assign   tb_o_ciphertext[887]                 =   tb_o_ciphertext[886];
assign   tb_o_tag_ready[887]                  =   1'b0;
assign   tb_o_tag[887]                        =   tb_o_tag[886];

// CLK no. 888/1240
// *************************************************
assign   tb_i_valid[888]                      =   1'b1;
assign   tb_i_reset[888]                      =   1'b0;
assign   tb_i_sop[888]                        =   1'b0;
assign   tb_i_key_update[888]                 =   1'b0;
assign   tb_i_key[888]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[888]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[888]               =   1'b0;
assign   tb_i_rf_static_encrypt[888]          =   1'b1;
assign   tb_i_clear_fault_flags[888]          =   1'b0;
assign   tb_i_rf_static_aad_length[888]       =   64'h0000000000000100;
assign   tb_i_aad[888]                        =   tb_i_aad[887];
assign   tb_i_rf_static_plaintext_length[888] =   64'h0000000000000280;
assign   tb_i_plaintext[888]                  =   256'h13e49006788c32756dcfa8cefc54b27fc1ce6050d28ddafc47b90b3f02287011;
assign   tb_o_valid[888]                      =   1'b0;
assign   tb_o_sop[888]                        =   1'b0;
assign   tb_o_ciphertext[888]                 =   tb_o_ciphertext[887];
assign   tb_o_tag_ready[888]                  =   1'b0;
assign   tb_o_tag[888]                        =   tb_o_tag[887];

// CLK no. 889/1240
// *************************************************
assign   tb_i_valid[889]                      =   1'b1;
assign   tb_i_reset[889]                      =   1'b0;
assign   tb_i_sop[889]                        =   1'b0;
assign   tb_i_key_update[889]                 =   1'b0;
assign   tb_i_key[889]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[889]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[889]               =   1'b0;
assign   tb_i_rf_static_encrypt[889]          =   1'b1;
assign   tb_i_clear_fault_flags[889]          =   1'b0;
assign   tb_i_rf_static_aad_length[889]       =   64'h0000000000000100;
assign   tb_i_aad[889]                        =   tb_i_aad[888];
assign   tb_i_rf_static_plaintext_length[889] =   64'h0000000000000280;
assign   tb_i_plaintext[889]                  =   256'hbeb6f65a53d592bb6aec28e2312ba1889422765c6e562584a51a9d158182fd3b;
assign   tb_o_valid[889]                      =   1'b0;
assign   tb_o_sop[889]                        =   1'b0;
assign   tb_o_ciphertext[889]                 =   tb_o_ciphertext[888];
assign   tb_o_tag_ready[889]                  =   1'b0;
assign   tb_o_tag[889]                        =   tb_o_tag[888];

// CLK no. 890/1240
// *************************************************
assign   tb_i_valid[890]                      =   1'b1;
assign   tb_i_reset[890]                      =   1'b0;
assign   tb_i_sop[890]                        =   1'b0;
assign   tb_i_key_update[890]                 =   1'b0;
assign   tb_i_key[890]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[890]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[890]               =   1'b0;
assign   tb_i_rf_static_encrypt[890]          =   1'b1;
assign   tb_i_clear_fault_flags[890]          =   1'b0;
assign   tb_i_rf_static_aad_length[890]       =   64'h0000000000000100;
assign   tb_i_aad[890]                        =   tb_i_aad[889];
assign   tb_i_rf_static_plaintext_length[890] =   64'h0000000000000280;
assign   tb_i_plaintext[890]                  =   256'h01e9d411754aa77afc6817e5c8ba0a07;
assign   tb_o_valid[890]                      =   1'b0;
assign   tb_o_sop[890]                        =   1'b0;
assign   tb_o_ciphertext[890]                 =   tb_o_ciphertext[889];
assign   tb_o_tag_ready[890]                  =   1'b0;
assign   tb_o_tag[890]                        =   tb_o_tag[889];

// CLK no. 891/1240
// *************************************************
assign   tb_i_valid[891]                      =   1'b0;
assign   tb_i_reset[891]                      =   1'b0;
assign   tb_i_sop[891]                        =   1'b0;
assign   tb_i_key_update[891]                 =   1'b0;
assign   tb_i_key[891]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[891]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[891]               =   1'b0;
assign   tb_i_rf_static_encrypt[891]          =   1'b1;
assign   tb_i_clear_fault_flags[891]          =   1'b0;
assign   tb_i_rf_static_aad_length[891]       =   64'h0000000000000100;
assign   tb_i_aad[891]                        =   tb_i_aad[890];
assign   tb_i_rf_static_plaintext_length[891] =   64'h0000000000000280;
assign   tb_i_plaintext[891]                  =   tb_i_plaintext[890];
assign   tb_o_valid[891]                      =   1'b0;
assign   tb_o_sop[891]                        =   1'b0;
assign   tb_o_ciphertext[891]                 =   tb_o_ciphertext[890];
assign   tb_o_tag_ready[891]                  =   1'b0;
assign   tb_o_tag[891]                        =   tb_o_tag[890];

// CLK no. 892/1240
// *************************************************
assign   tb_i_valid[892]                      =   1'b0;
assign   tb_i_reset[892]                      =   1'b0;
assign   tb_i_sop[892]                        =   1'b0;
assign   tb_i_key_update[892]                 =   1'b0;
assign   tb_i_key[892]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[892]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[892]               =   1'b0;
assign   tb_i_rf_static_encrypt[892]          =   1'b1;
assign   tb_i_clear_fault_flags[892]          =   1'b0;
assign   tb_i_rf_static_aad_length[892]       =   64'h0000000000000100;
assign   tb_i_aad[892]                        =   tb_i_aad[891];
assign   tb_i_rf_static_plaintext_length[892] =   64'h0000000000000280;
assign   tb_i_plaintext[892]                  =   tb_i_plaintext[891];
assign   tb_o_valid[892]                      =   1'b0;
assign   tb_o_sop[892]                        =   1'b0;
assign   tb_o_ciphertext[892]                 =   tb_o_ciphertext[891];
assign   tb_o_tag_ready[892]                  =   1'b0;
assign   tb_o_tag[892]                        =   tb_o_tag[891];

// CLK no. 893/1240
// *************************************************
assign   tb_i_valid[893]                      =   1'b0;
assign   tb_i_reset[893]                      =   1'b0;
assign   tb_i_sop[893]                        =   1'b0;
assign   tb_i_key_update[893]                 =   1'b0;
assign   tb_i_key[893]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[893]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[893]               =   1'b0;
assign   tb_i_rf_static_encrypt[893]          =   1'b1;
assign   tb_i_clear_fault_flags[893]          =   1'b0;
assign   tb_i_rf_static_aad_length[893]       =   64'h0000000000000100;
assign   tb_i_aad[893]                        =   tb_i_aad[892];
assign   tb_i_rf_static_plaintext_length[893] =   64'h0000000000000280;
assign   tb_i_plaintext[893]                  =   tb_i_plaintext[892];
assign   tb_o_valid[893]                      =   1'b0;
assign   tb_o_sop[893]                        =   1'b0;
assign   tb_o_ciphertext[893]                 =   tb_o_ciphertext[892];
assign   tb_o_tag_ready[893]                  =   1'b0;
assign   tb_o_tag[893]                        =   tb_o_tag[892];

// CLK no. 894/1240
// *************************************************
assign   tb_i_valid[894]                      =   1'b0;
assign   tb_i_reset[894]                      =   1'b0;
assign   tb_i_sop[894]                        =   1'b0;
assign   tb_i_key_update[894]                 =   1'b0;
assign   tb_i_key[894]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[894]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[894]               =   1'b0;
assign   tb_i_rf_static_encrypt[894]          =   1'b1;
assign   tb_i_clear_fault_flags[894]          =   1'b0;
assign   tb_i_rf_static_aad_length[894]       =   64'h0000000000000100;
assign   tb_i_aad[894]                        =   tb_i_aad[893];
assign   tb_i_rf_static_plaintext_length[894] =   64'h0000000000000280;
assign   tb_i_plaintext[894]                  =   tb_i_plaintext[893];
assign   tb_o_valid[894]                      =   1'b0;
assign   tb_o_sop[894]                        =   1'b0;
assign   tb_o_ciphertext[894]                 =   tb_o_ciphertext[893];
assign   tb_o_tag_ready[894]                  =   1'b0;
assign   tb_o_tag[894]                        =   tb_o_tag[893];

// CLK no. 895/1240
// *************************************************
assign   tb_i_valid[895]                      =   1'b0;
assign   tb_i_reset[895]                      =   1'b0;
assign   tb_i_sop[895]                        =   1'b0;
assign   tb_i_key_update[895]                 =   1'b0;
assign   tb_i_key[895]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[895]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[895]               =   1'b0;
assign   tb_i_rf_static_encrypt[895]          =   1'b1;
assign   tb_i_clear_fault_flags[895]          =   1'b0;
assign   tb_i_rf_static_aad_length[895]       =   64'h0000000000000100;
assign   tb_i_aad[895]                        =   tb_i_aad[894];
assign   tb_i_rf_static_plaintext_length[895] =   64'h0000000000000280;
assign   tb_i_plaintext[895]                  =   tb_i_plaintext[894];
assign   tb_o_valid[895]                      =   1'b0;
assign   tb_o_sop[895]                        =   1'b0;
assign   tb_o_ciphertext[895]                 =   tb_o_ciphertext[894];
assign   tb_o_tag_ready[895]                  =   1'b0;
assign   tb_o_tag[895]                        =   tb_o_tag[894];

// CLK no. 896/1240
// *************************************************
assign   tb_i_valid[896]                      =   1'b0;
assign   tb_i_reset[896]                      =   1'b0;
assign   tb_i_sop[896]                        =   1'b0;
assign   tb_i_key_update[896]                 =   1'b0;
assign   tb_i_key[896]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[896]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[896]               =   1'b0;
assign   tb_i_rf_static_encrypt[896]          =   1'b1;
assign   tb_i_clear_fault_flags[896]          =   1'b0;
assign   tb_i_rf_static_aad_length[896]       =   64'h0000000000000100;
assign   tb_i_aad[896]                        =   tb_i_aad[895];
assign   tb_i_rf_static_plaintext_length[896] =   64'h0000000000000280;
assign   tb_i_plaintext[896]                  =   tb_i_plaintext[895];
assign   tb_o_valid[896]                      =   1'b0;
assign   tb_o_sop[896]                        =   1'b0;
assign   tb_o_ciphertext[896]                 =   tb_o_ciphertext[895];
assign   tb_o_tag_ready[896]                  =   1'b0;
assign   tb_o_tag[896]                        =   tb_o_tag[895];

// CLK no. 897/1240
// *************************************************
assign   tb_i_valid[897]                      =   1'b0;
assign   tb_i_reset[897]                      =   1'b0;
assign   tb_i_sop[897]                        =   1'b0;
assign   tb_i_key_update[897]                 =   1'b0;
assign   tb_i_key[897]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[897]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[897]               =   1'b0;
assign   tb_i_rf_static_encrypt[897]          =   1'b1;
assign   tb_i_clear_fault_flags[897]          =   1'b0;
assign   tb_i_rf_static_aad_length[897]       =   64'h0000000000000100;
assign   tb_i_aad[897]                        =   tb_i_aad[896];
assign   tb_i_rf_static_plaintext_length[897] =   64'h0000000000000280;
assign   tb_i_plaintext[897]                  =   tb_i_plaintext[896];
assign   tb_o_valid[897]                      =   1'b0;
assign   tb_o_sop[897]                        =   1'b0;
assign   tb_o_ciphertext[897]                 =   tb_o_ciphertext[896];
assign   tb_o_tag_ready[897]                  =   1'b0;
assign   tb_o_tag[897]                        =   tb_o_tag[896];

// CLK no. 898/1240
// *************************************************
assign   tb_i_valid[898]                      =   1'b0;
assign   tb_i_reset[898]                      =   1'b0;
assign   tb_i_sop[898]                        =   1'b0;
assign   tb_i_key_update[898]                 =   1'b0;
assign   tb_i_key[898]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[898]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[898]               =   1'b0;
assign   tb_i_rf_static_encrypt[898]          =   1'b1;
assign   tb_i_clear_fault_flags[898]          =   1'b0;
assign   tb_i_rf_static_aad_length[898]       =   64'h0000000000000100;
assign   tb_i_aad[898]                        =   tb_i_aad[897];
assign   tb_i_rf_static_plaintext_length[898] =   64'h0000000000000280;
assign   tb_i_plaintext[898]                  =   tb_i_plaintext[897];
assign   tb_o_valid[898]                      =   1'b0;
assign   tb_o_sop[898]                        =   1'b0;
assign   tb_o_ciphertext[898]                 =   tb_o_ciphertext[897];
assign   tb_o_tag_ready[898]                  =   1'b0;
assign   tb_o_tag[898]                        =   tb_o_tag[897];

// CLK no. 899/1240
// *************************************************
assign   tb_i_valid[899]                      =   1'b0;
assign   tb_i_reset[899]                      =   1'b0;
assign   tb_i_sop[899]                        =   1'b0;
assign   tb_i_key_update[899]                 =   1'b0;
assign   tb_i_key[899]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[899]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[899]               =   1'b0;
assign   tb_i_rf_static_encrypt[899]          =   1'b1;
assign   tb_i_clear_fault_flags[899]          =   1'b0;
assign   tb_i_rf_static_aad_length[899]       =   64'h0000000000000100;
assign   tb_i_aad[899]                        =   tb_i_aad[898];
assign   tb_i_rf_static_plaintext_length[899] =   64'h0000000000000280;
assign   tb_i_plaintext[899]                  =   tb_i_plaintext[898];
assign   tb_o_valid[899]                      =   1'b0;
assign   tb_o_sop[899]                        =   1'b0;
assign   tb_o_ciphertext[899]                 =   tb_o_ciphertext[898];
assign   tb_o_tag_ready[899]                  =   1'b0;
assign   tb_o_tag[899]                        =   tb_o_tag[898];

// CLK no. 900/1240
// *************************************************
assign   tb_i_valid[900]                      =   1'b0;
assign   tb_i_reset[900]                      =   1'b0;
assign   tb_i_sop[900]                        =   1'b0;
assign   tb_i_key_update[900]                 =   1'b0;
assign   tb_i_key[900]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[900]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[900]               =   1'b0;
assign   tb_i_rf_static_encrypt[900]          =   1'b1;
assign   tb_i_clear_fault_flags[900]          =   1'b0;
assign   tb_i_rf_static_aad_length[900]       =   64'h0000000000000100;
assign   tb_i_aad[900]                        =   tb_i_aad[899];
assign   tb_i_rf_static_plaintext_length[900] =   64'h0000000000000280;
assign   tb_i_plaintext[900]                  =   tb_i_plaintext[899];
assign   tb_o_valid[900]                      =   1'b0;
assign   tb_o_sop[900]                        =   1'b0;
assign   tb_o_ciphertext[900]                 =   tb_o_ciphertext[899];
assign   tb_o_tag_ready[900]                  =   1'b0;
assign   tb_o_tag[900]                        =   tb_o_tag[899];

// CLK no. 901/1240
// *************************************************
assign   tb_i_valid[901]                      =   1'b0;
assign   tb_i_reset[901]                      =   1'b0;
assign   tb_i_sop[901]                        =   1'b0;
assign   tb_i_key_update[901]                 =   1'b0;
assign   tb_i_key[901]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[901]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[901]               =   1'b0;
assign   tb_i_rf_static_encrypt[901]          =   1'b1;
assign   tb_i_clear_fault_flags[901]          =   1'b0;
assign   tb_i_rf_static_aad_length[901]       =   64'h0000000000000100;
assign   tb_i_aad[901]                        =   tb_i_aad[900];
assign   tb_i_rf_static_plaintext_length[901] =   64'h0000000000000280;
assign   tb_i_plaintext[901]                  =   tb_i_plaintext[900];
assign   tb_o_valid[901]                      =   1'b0;
assign   tb_o_sop[901]                        =   1'b0;
assign   tb_o_ciphertext[901]                 =   tb_o_ciphertext[900];
assign   tb_o_tag_ready[901]                  =   1'b0;
assign   tb_o_tag[901]                        =   tb_o_tag[900];

// CLK no. 902/1240
// *************************************************
assign   tb_i_valid[902]                      =   1'b0;
assign   tb_i_reset[902]                      =   1'b0;
assign   tb_i_sop[902]                        =   1'b0;
assign   tb_i_key_update[902]                 =   1'b0;
assign   tb_i_key[902]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[902]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[902]               =   1'b0;
assign   tb_i_rf_static_encrypt[902]          =   1'b1;
assign   tb_i_clear_fault_flags[902]          =   1'b0;
assign   tb_i_rf_static_aad_length[902]       =   64'h0000000000000100;
assign   tb_i_aad[902]                        =   tb_i_aad[901];
assign   tb_i_rf_static_plaintext_length[902] =   64'h0000000000000280;
assign   tb_i_plaintext[902]                  =   tb_i_plaintext[901];
assign   tb_o_valid[902]                      =   1'b0;
assign   tb_o_sop[902]                        =   1'b0;
assign   tb_o_ciphertext[902]                 =   tb_o_ciphertext[901];
assign   tb_o_tag_ready[902]                  =   1'b0;
assign   tb_o_tag[902]                        =   tb_o_tag[901];

// CLK no. 903/1240
// *************************************************
assign   tb_i_valid[903]                      =   1'b0;
assign   tb_i_reset[903]                      =   1'b0;
assign   tb_i_sop[903]                        =   1'b0;
assign   tb_i_key_update[903]                 =   1'b0;
assign   tb_i_key[903]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[903]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[903]               =   1'b0;
assign   tb_i_rf_static_encrypt[903]          =   1'b1;
assign   tb_i_clear_fault_flags[903]          =   1'b0;
assign   tb_i_rf_static_aad_length[903]       =   64'h0000000000000100;
assign   tb_i_aad[903]                        =   tb_i_aad[902];
assign   tb_i_rf_static_plaintext_length[903] =   64'h0000000000000280;
assign   tb_i_plaintext[903]                  =   tb_i_plaintext[902];
assign   tb_o_valid[903]                      =   1'b0;
assign   tb_o_sop[903]                        =   1'b0;
assign   tb_o_ciphertext[903]                 =   tb_o_ciphertext[902];
assign   tb_o_tag_ready[903]                  =   1'b0;
assign   tb_o_tag[903]                        =   tb_o_tag[902];

// CLK no. 904/1240
// *************************************************
assign   tb_i_valid[904]                      =   1'b0;
assign   tb_i_reset[904]                      =   1'b0;
assign   tb_i_sop[904]                        =   1'b0;
assign   tb_i_key_update[904]                 =   1'b0;
assign   tb_i_key[904]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[904]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[904]               =   1'b0;
assign   tb_i_rf_static_encrypt[904]          =   1'b1;
assign   tb_i_clear_fault_flags[904]          =   1'b0;
assign   tb_i_rf_static_aad_length[904]       =   64'h0000000000000100;
assign   tb_i_aad[904]                        =   tb_i_aad[903];
assign   tb_i_rf_static_plaintext_length[904] =   64'h0000000000000280;
assign   tb_i_plaintext[904]                  =   tb_i_plaintext[903];
assign   tb_o_valid[904]                      =   1'b0;
assign   tb_o_sop[904]                        =   1'b0;
assign   tb_o_ciphertext[904]                 =   tb_o_ciphertext[903];
assign   tb_o_tag_ready[904]                  =   1'b0;
assign   tb_o_tag[904]                        =   tb_o_tag[903];

// CLK no. 905/1240
// *************************************************
assign   tb_i_valid[905]                      =   1'b0;
assign   tb_i_reset[905]                      =   1'b0;
assign   tb_i_sop[905]                        =   1'b0;
assign   tb_i_key_update[905]                 =   1'b0;
assign   tb_i_key[905]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[905]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[905]               =   1'b0;
assign   tb_i_rf_static_encrypt[905]          =   1'b1;
assign   tb_i_clear_fault_flags[905]          =   1'b0;
assign   tb_i_rf_static_aad_length[905]       =   64'h0000000000000100;
assign   tb_i_aad[905]                        =   tb_i_aad[904];
assign   tb_i_rf_static_plaintext_length[905] =   64'h0000000000000280;
assign   tb_i_plaintext[905]                  =   tb_i_plaintext[904];
assign   tb_o_valid[905]                      =   1'b0;
assign   tb_o_sop[905]                        =   1'b0;
assign   tb_o_ciphertext[905]                 =   tb_o_ciphertext[904];
assign   tb_o_tag_ready[905]                  =   1'b0;
assign   tb_o_tag[905]                        =   tb_o_tag[904];

// CLK no. 906/1240
// *************************************************
assign   tb_i_valid[906]                      =   1'b0;
assign   tb_i_reset[906]                      =   1'b0;
assign   tb_i_sop[906]                        =   1'b0;
assign   tb_i_key_update[906]                 =   1'b0;
assign   tb_i_key[906]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[906]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[906]               =   1'b0;
assign   tb_i_rf_static_encrypt[906]          =   1'b1;
assign   tb_i_clear_fault_flags[906]          =   1'b0;
assign   tb_i_rf_static_aad_length[906]       =   64'h0000000000000100;
assign   tb_i_aad[906]                        =   tb_i_aad[905];
assign   tb_i_rf_static_plaintext_length[906] =   64'h0000000000000280;
assign   tb_i_plaintext[906]                  =   tb_i_plaintext[905];
assign   tb_o_valid[906]                      =   1'b0;
assign   tb_o_sop[906]                        =   1'b0;
assign   tb_o_ciphertext[906]                 =   tb_o_ciphertext[905];
assign   tb_o_tag_ready[906]                  =   1'b0;
assign   tb_o_tag[906]                        =   tb_o_tag[905];

// CLK no. 907/1240
// *************************************************
assign   tb_i_valid[907]                      =   1'b0;
assign   tb_i_reset[907]                      =   1'b0;
assign   tb_i_sop[907]                        =   1'b0;
assign   tb_i_key_update[907]                 =   1'b0;
assign   tb_i_key[907]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[907]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[907]               =   1'b0;
assign   tb_i_rf_static_encrypt[907]          =   1'b1;
assign   tb_i_clear_fault_flags[907]          =   1'b0;
assign   tb_i_rf_static_aad_length[907]       =   64'h0000000000000100;
assign   tb_i_aad[907]                        =   tb_i_aad[906];
assign   tb_i_rf_static_plaintext_length[907] =   64'h0000000000000280;
assign   tb_i_plaintext[907]                  =   tb_i_plaintext[906];
assign   tb_o_valid[907]                      =   1'b0;
assign   tb_o_sop[907]                        =   1'b0;
assign   tb_o_ciphertext[907]                 =   tb_o_ciphertext[906];
assign   tb_o_tag_ready[907]                  =   1'b0;
assign   tb_o_tag[907]                        =   tb_o_tag[906];

// CLK no. 908/1240
// *************************************************
assign   tb_i_valid[908]                      =   1'b0;
assign   tb_i_reset[908]                      =   1'b0;
assign   tb_i_sop[908]                        =   1'b0;
assign   tb_i_key_update[908]                 =   1'b0;
assign   tb_i_key[908]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[908]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[908]               =   1'b0;
assign   tb_i_rf_static_encrypt[908]          =   1'b1;
assign   tb_i_clear_fault_flags[908]          =   1'b0;
assign   tb_i_rf_static_aad_length[908]       =   64'h0000000000000100;
assign   tb_i_aad[908]                        =   tb_i_aad[907];
assign   tb_i_rf_static_plaintext_length[908] =   64'h0000000000000280;
assign   tb_i_plaintext[908]                  =   tb_i_plaintext[907];
assign   tb_o_valid[908]                      =   1'b0;
assign   tb_o_sop[908]                        =   1'b0;
assign   tb_o_ciphertext[908]                 =   tb_o_ciphertext[907];
assign   tb_o_tag_ready[908]                  =   1'b0;
assign   tb_o_tag[908]                        =   tb_o_tag[907];

// CLK no. 909/1240
// *************************************************
assign   tb_i_valid[909]                      =   1'b0;
assign   tb_i_reset[909]                      =   1'b0;
assign   tb_i_sop[909]                        =   1'b0;
assign   tb_i_key_update[909]                 =   1'b0;
assign   tb_i_key[909]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[909]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[909]               =   1'b0;
assign   tb_i_rf_static_encrypt[909]          =   1'b1;
assign   tb_i_clear_fault_flags[909]          =   1'b0;
assign   tb_i_rf_static_aad_length[909]       =   64'h0000000000000100;
assign   tb_i_aad[909]                        =   tb_i_aad[908];
assign   tb_i_rf_static_plaintext_length[909] =   64'h0000000000000280;
assign   tb_i_plaintext[909]                  =   tb_i_plaintext[908];
assign   tb_o_valid[909]                      =   1'b0;
assign   tb_o_sop[909]                        =   1'b0;
assign   tb_o_ciphertext[909]                 =   tb_o_ciphertext[908];
assign   tb_o_tag_ready[909]                  =   1'b0;
assign   tb_o_tag[909]                        =   tb_o_tag[908];

// CLK no. 910/1240
// *************************************************
assign   tb_i_valid[910]                      =   1'b0;
assign   tb_i_reset[910]                      =   1'b0;
assign   tb_i_sop[910]                        =   1'b0;
assign   tb_i_key_update[910]                 =   1'b0;
assign   tb_i_key[910]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[910]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[910]               =   1'b0;
assign   tb_i_rf_static_encrypt[910]          =   1'b1;
assign   tb_i_clear_fault_flags[910]          =   1'b0;
assign   tb_i_rf_static_aad_length[910]       =   64'h0000000000000100;
assign   tb_i_aad[910]                        =   tb_i_aad[909];
assign   tb_i_rf_static_plaintext_length[910] =   64'h0000000000000280;
assign   tb_i_plaintext[910]                  =   tb_i_plaintext[909];
assign   tb_o_valid[910]                      =   1'b0;
assign   tb_o_sop[910]                        =   1'b0;
assign   tb_o_ciphertext[910]                 =   tb_o_ciphertext[909];
assign   tb_o_tag_ready[910]                  =   1'b0;
assign   tb_o_tag[910]                        =   tb_o_tag[909];

// CLK no. 911/1240
// *************************************************
assign   tb_i_valid[911]                      =   1'b0;
assign   tb_i_reset[911]                      =   1'b0;
assign   tb_i_sop[911]                        =   1'b0;
assign   tb_i_key_update[911]                 =   1'b0;
assign   tb_i_key[911]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[911]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[911]               =   1'b0;
assign   tb_i_rf_static_encrypt[911]          =   1'b1;
assign   tb_i_clear_fault_flags[911]          =   1'b0;
assign   tb_i_rf_static_aad_length[911]       =   64'h0000000000000100;
assign   tb_i_aad[911]                        =   tb_i_aad[910];
assign   tb_i_rf_static_plaintext_length[911] =   64'h0000000000000280;
assign   tb_i_plaintext[911]                  =   tb_i_plaintext[910];
assign   tb_o_valid[911]                      =   1'b0;
assign   tb_o_sop[911]                        =   1'b0;
assign   tb_o_ciphertext[911]                 =   tb_o_ciphertext[910];
assign   tb_o_tag_ready[911]                  =   1'b0;
assign   tb_o_tag[911]                        =   tb_o_tag[910];

// CLK no. 912/1240
// *************************************************
assign   tb_i_valid[912]                      =   1'b0;
assign   tb_i_reset[912]                      =   1'b0;
assign   tb_i_sop[912]                        =   1'b0;
assign   tb_i_key_update[912]                 =   1'b0;
assign   tb_i_key[912]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[912]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[912]               =   1'b0;
assign   tb_i_rf_static_encrypt[912]          =   1'b1;
assign   tb_i_clear_fault_flags[912]          =   1'b0;
assign   tb_i_rf_static_aad_length[912]       =   64'h0000000000000100;
assign   tb_i_aad[912]                        =   tb_i_aad[911];
assign   tb_i_rf_static_plaintext_length[912] =   64'h0000000000000280;
assign   tb_i_plaintext[912]                  =   tb_i_plaintext[911];
assign   tb_o_valid[912]                      =   1'b0;
assign   tb_o_sop[912]                        =   1'b0;
assign   tb_o_ciphertext[912]                 =   tb_o_ciphertext[911];
assign   tb_o_tag_ready[912]                  =   1'b0;
assign   tb_o_tag[912]                        =   tb_o_tag[911];

// CLK no. 913/1240
// *************************************************
assign   tb_i_valid[913]                      =   1'b0;
assign   tb_i_reset[913]                      =   1'b0;
assign   tb_i_sop[913]                        =   1'b0;
assign   tb_i_key_update[913]                 =   1'b0;
assign   tb_i_key[913]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[913]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[913]               =   1'b0;
assign   tb_i_rf_static_encrypt[913]          =   1'b1;
assign   tb_i_clear_fault_flags[913]          =   1'b0;
assign   tb_i_rf_static_aad_length[913]       =   64'h0000000000000100;
assign   tb_i_aad[913]                        =   tb_i_aad[912];
assign   tb_i_rf_static_plaintext_length[913] =   64'h0000000000000280;
assign   tb_i_plaintext[913]                  =   tb_i_plaintext[912];
assign   tb_o_valid[913]                      =   1'b0;
assign   tb_o_sop[913]                        =   1'b0;
assign   tb_o_ciphertext[913]                 =   tb_o_ciphertext[912];
assign   tb_o_tag_ready[913]                  =   1'b0;
assign   tb_o_tag[913]                        =   tb_o_tag[912];

// CLK no. 914/1240
// *************************************************
assign   tb_i_valid[914]                      =   1'b0;
assign   tb_i_reset[914]                      =   1'b0;
assign   tb_i_sop[914]                        =   1'b0;
assign   tb_i_key_update[914]                 =   1'b0;
assign   tb_i_key[914]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[914]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[914]               =   1'b0;
assign   tb_i_rf_static_encrypt[914]          =   1'b1;
assign   tb_i_clear_fault_flags[914]          =   1'b0;
assign   tb_i_rf_static_aad_length[914]       =   64'h0000000000000100;
assign   tb_i_aad[914]                        =   tb_i_aad[913];
assign   tb_i_rf_static_plaintext_length[914] =   64'h0000000000000280;
assign   tb_i_plaintext[914]                  =   tb_i_plaintext[913];
assign   tb_o_valid[914]                      =   1'b0;
assign   tb_o_sop[914]                        =   1'b0;
assign   tb_o_ciphertext[914]                 =   tb_o_ciphertext[913];
assign   tb_o_tag_ready[914]                  =   1'b0;
assign   tb_o_tag[914]                        =   tb_o_tag[913];

// CLK no. 915/1240
// *************************************************
assign   tb_i_valid[915]                      =   1'b0;
assign   tb_i_reset[915]                      =   1'b0;
assign   tb_i_sop[915]                        =   1'b0;
assign   tb_i_key_update[915]                 =   1'b0;
assign   tb_i_key[915]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[915]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[915]               =   1'b0;
assign   tb_i_rf_static_encrypt[915]          =   1'b1;
assign   tb_i_clear_fault_flags[915]          =   1'b0;
assign   tb_i_rf_static_aad_length[915]       =   64'h0000000000000100;
assign   tb_i_aad[915]                        =   tb_i_aad[914];
assign   tb_i_rf_static_plaintext_length[915] =   64'h0000000000000280;
assign   tb_i_plaintext[915]                  =   tb_i_plaintext[914];
assign   tb_o_valid[915]                      =   1'b0;
assign   tb_o_sop[915]                        =   1'b0;
assign   tb_o_ciphertext[915]                 =   tb_o_ciphertext[914];
assign   tb_o_tag_ready[915]                  =   1'b0;
assign   tb_o_tag[915]                        =   tb_o_tag[914];

// CLK no. 916/1240
// *************************************************
assign   tb_i_valid[916]                      =   1'b0;
assign   tb_i_reset[916]                      =   1'b0;
assign   tb_i_sop[916]                        =   1'b0;
assign   tb_i_key_update[916]                 =   1'b0;
assign   tb_i_key[916]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[916]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[916]               =   1'b0;
assign   tb_i_rf_static_encrypt[916]          =   1'b1;
assign   tb_i_clear_fault_flags[916]          =   1'b0;
assign   tb_i_rf_static_aad_length[916]       =   64'h0000000000000100;
assign   tb_i_aad[916]                        =   tb_i_aad[915];
assign   tb_i_rf_static_plaintext_length[916] =   64'h0000000000000280;
assign   tb_i_plaintext[916]                  =   tb_i_plaintext[915];
assign   tb_o_valid[916]                      =   1'b0;
assign   tb_o_sop[916]                        =   1'b0;
assign   tb_o_ciphertext[916]                 =   tb_o_ciphertext[915];
assign   tb_o_tag_ready[916]                  =   1'b0;
assign   tb_o_tag[916]                        =   tb_o_tag[915];

// CLK no. 917/1240
// *************************************************
assign   tb_i_valid[917]                      =   1'b0;
assign   tb_i_reset[917]                      =   1'b0;
assign   tb_i_sop[917]                        =   1'b0;
assign   tb_i_key_update[917]                 =   1'b0;
assign   tb_i_key[917]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[917]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[917]               =   1'b0;
assign   tb_i_rf_static_encrypt[917]          =   1'b1;
assign   tb_i_clear_fault_flags[917]          =   1'b0;
assign   tb_i_rf_static_aad_length[917]       =   64'h0000000000000100;
assign   tb_i_aad[917]                        =   tb_i_aad[916];
assign   tb_i_rf_static_plaintext_length[917] =   64'h0000000000000280;
assign   tb_i_plaintext[917]                  =   tb_i_plaintext[916];
assign   tb_o_valid[917]                      =   1'b0;
assign   tb_o_sop[917]                        =   1'b0;
assign   tb_o_ciphertext[917]                 =   tb_o_ciphertext[916];
assign   tb_o_tag_ready[917]                  =   1'b0;
assign   tb_o_tag[917]                        =   tb_o_tag[916];

// CLK no. 918/1240
// *************************************************
assign   tb_i_valid[918]                      =   1'b0;
assign   tb_i_reset[918]                      =   1'b0;
assign   tb_i_sop[918]                        =   1'b0;
assign   tb_i_key_update[918]                 =   1'b0;
assign   tb_i_key[918]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[918]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[918]               =   1'b0;
assign   tb_i_rf_static_encrypt[918]          =   1'b1;
assign   tb_i_clear_fault_flags[918]          =   1'b0;
assign   tb_i_rf_static_aad_length[918]       =   64'h0000000000000100;
assign   tb_i_aad[918]                        =   tb_i_aad[917];
assign   tb_i_rf_static_plaintext_length[918] =   64'h0000000000000280;
assign   tb_i_plaintext[918]                  =   tb_i_plaintext[917];
assign   tb_o_valid[918]                      =   1'b0;
assign   tb_o_sop[918]                        =   1'b0;
assign   tb_o_ciphertext[918]                 =   tb_o_ciphertext[917];
assign   tb_o_tag_ready[918]                  =   1'b0;
assign   tb_o_tag[918]                        =   tb_o_tag[917];

// CLK no. 919/1240
// *************************************************
assign   tb_i_valid[919]                      =   1'b0;
assign   tb_i_reset[919]                      =   1'b0;
assign   tb_i_sop[919]                        =   1'b0;
assign   tb_i_key_update[919]                 =   1'b0;
assign   tb_i_key[919]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[919]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[919]               =   1'b0;
assign   tb_i_rf_static_encrypt[919]          =   1'b1;
assign   tb_i_clear_fault_flags[919]          =   1'b0;
assign   tb_i_rf_static_aad_length[919]       =   64'h0000000000000100;
assign   tb_i_aad[919]                        =   tb_i_aad[918];
assign   tb_i_rf_static_plaintext_length[919] =   64'h0000000000000280;
assign   tb_i_plaintext[919]                  =   tb_i_plaintext[918];
assign   tb_o_valid[919]                      =   1'b0;
assign   tb_o_sop[919]                        =   1'b0;
assign   tb_o_ciphertext[919]                 =   tb_o_ciphertext[918];
assign   tb_o_tag_ready[919]                  =   1'b0;
assign   tb_o_tag[919]                        =   tb_o_tag[918];

// CLK no. 920/1240
// *************************************************
assign   tb_i_valid[920]                      =   1'b0;
assign   tb_i_reset[920]                      =   1'b0;
assign   tb_i_sop[920]                        =   1'b0;
assign   tb_i_key_update[920]                 =   1'b0;
assign   tb_i_key[920]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[920]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[920]               =   1'b0;
assign   tb_i_rf_static_encrypt[920]          =   1'b1;
assign   tb_i_clear_fault_flags[920]          =   1'b0;
assign   tb_i_rf_static_aad_length[920]       =   64'h0000000000000100;
assign   tb_i_aad[920]                        =   tb_i_aad[919];
assign   tb_i_rf_static_plaintext_length[920] =   64'h0000000000000280;
assign   tb_i_plaintext[920]                  =   tb_i_plaintext[919];
assign   tb_o_valid[920]                      =   1'b0;
assign   tb_o_sop[920]                        =   1'b0;
assign   tb_o_ciphertext[920]                 =   tb_o_ciphertext[919];
assign   tb_o_tag_ready[920]                  =   1'b0;
assign   tb_o_tag[920]                        =   tb_o_tag[919];

// CLK no. 921/1240
// *************************************************
assign   tb_i_valid[921]                      =   1'b0;
assign   tb_i_reset[921]                      =   1'b0;
assign   tb_i_sop[921]                        =   1'b0;
assign   tb_i_key_update[921]                 =   1'b0;
assign   tb_i_key[921]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[921]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[921]               =   1'b0;
assign   tb_i_rf_static_encrypt[921]          =   1'b1;
assign   tb_i_clear_fault_flags[921]          =   1'b0;
assign   tb_i_rf_static_aad_length[921]       =   64'h0000000000000100;
assign   tb_i_aad[921]                        =   tb_i_aad[920];
assign   tb_i_rf_static_plaintext_length[921] =   64'h0000000000000280;
assign   tb_i_plaintext[921]                  =   tb_i_plaintext[920];
assign   tb_o_valid[921]                      =   1'b0;
assign   tb_o_sop[921]                        =   1'b0;
assign   tb_o_ciphertext[921]                 =   tb_o_ciphertext[920];
assign   tb_o_tag_ready[921]                  =   1'b0;
assign   tb_o_tag[921]                        =   tb_o_tag[920];

// CLK no. 922/1240
// *************************************************
assign   tb_i_valid[922]                      =   1'b0;
assign   tb_i_reset[922]                      =   1'b0;
assign   tb_i_sop[922]                        =   1'b0;
assign   tb_i_key_update[922]                 =   1'b0;
assign   tb_i_key[922]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[922]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[922]               =   1'b0;
assign   tb_i_rf_static_encrypt[922]          =   1'b1;
assign   tb_i_clear_fault_flags[922]          =   1'b0;
assign   tb_i_rf_static_aad_length[922]       =   64'h0000000000000100;
assign   tb_i_aad[922]                        =   tb_i_aad[921];
assign   tb_i_rf_static_plaintext_length[922] =   64'h0000000000000280;
assign   tb_i_plaintext[922]                  =   tb_i_plaintext[921];
assign   tb_o_valid[922]                      =   1'b0;
assign   tb_o_sop[922]                        =   1'b0;
assign   tb_o_ciphertext[922]                 =   tb_o_ciphertext[921];
assign   tb_o_tag_ready[922]                  =   1'b0;
assign   tb_o_tag[922]                        =   tb_o_tag[921];

// CLK no. 923/1240
// *************************************************
assign   tb_i_valid[923]                      =   1'b0;
assign   tb_i_reset[923]                      =   1'b0;
assign   tb_i_sop[923]                        =   1'b0;
assign   tb_i_key_update[923]                 =   1'b0;
assign   tb_i_key[923]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[923]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[923]               =   1'b0;
assign   tb_i_rf_static_encrypt[923]          =   1'b1;
assign   tb_i_clear_fault_flags[923]          =   1'b0;
assign   tb_i_rf_static_aad_length[923]       =   64'h0000000000000100;
assign   tb_i_aad[923]                        =   tb_i_aad[922];
assign   tb_i_rf_static_plaintext_length[923] =   64'h0000000000000280;
assign   tb_i_plaintext[923]                  =   tb_i_plaintext[922];
assign   tb_o_valid[923]                      =   1'b0;
assign   tb_o_sop[923]                        =   1'b0;
assign   tb_o_ciphertext[923]                 =   tb_o_ciphertext[922];
assign   tb_o_tag_ready[923]                  =   1'b0;
assign   tb_o_tag[923]                        =   tb_o_tag[922];

// CLK no. 924/1240
// *************************************************
assign   tb_i_valid[924]                      =   1'b0;
assign   tb_i_reset[924]                      =   1'b0;
assign   tb_i_sop[924]                        =   1'b0;
assign   tb_i_key_update[924]                 =   1'b0;
assign   tb_i_key[924]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[924]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[924]               =   1'b0;
assign   tb_i_rf_static_encrypt[924]          =   1'b1;
assign   tb_i_clear_fault_flags[924]          =   1'b0;
assign   tb_i_rf_static_aad_length[924]       =   64'h0000000000000100;
assign   tb_i_aad[924]                        =   tb_i_aad[923];
assign   tb_i_rf_static_plaintext_length[924] =   64'h0000000000000280;
assign   tb_i_plaintext[924]                  =   tb_i_plaintext[923];
assign   tb_o_valid[924]                      =   1'b0;
assign   tb_o_sop[924]                        =   1'b0;
assign   tb_o_ciphertext[924]                 =   tb_o_ciphertext[923];
assign   tb_o_tag_ready[924]                  =   1'b0;
assign   tb_o_tag[924]                        =   tb_o_tag[923];

// CLK no. 925/1240
// *************************************************
assign   tb_i_valid[925]                      =   1'b0;
assign   tb_i_reset[925]                      =   1'b0;
assign   tb_i_sop[925]                        =   1'b0;
assign   tb_i_key_update[925]                 =   1'b0;
assign   tb_i_key[925]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[925]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[925]               =   1'b0;
assign   tb_i_rf_static_encrypt[925]          =   1'b1;
assign   tb_i_clear_fault_flags[925]          =   1'b0;
assign   tb_i_rf_static_aad_length[925]       =   64'h0000000000000100;
assign   tb_i_aad[925]                        =   tb_i_aad[924];
assign   tb_i_rf_static_plaintext_length[925] =   64'h0000000000000280;
assign   tb_i_plaintext[925]                  =   tb_i_plaintext[924];
assign   tb_o_valid[925]                      =   1'b0;
assign   tb_o_sop[925]                        =   1'b0;
assign   tb_o_ciphertext[925]                 =   tb_o_ciphertext[924];
assign   tb_o_tag_ready[925]                  =   1'b0;
assign   tb_o_tag[925]                        =   tb_o_tag[924];

// CLK no. 926/1240
// *************************************************
assign   tb_i_valid[926]                      =   1'b0;
assign   tb_i_reset[926]                      =   1'b0;
assign   tb_i_sop[926]                        =   1'b0;
assign   tb_i_key_update[926]                 =   1'b0;
assign   tb_i_key[926]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[926]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[926]               =   1'b0;
assign   tb_i_rf_static_encrypt[926]          =   1'b1;
assign   tb_i_clear_fault_flags[926]          =   1'b0;
assign   tb_i_rf_static_aad_length[926]       =   64'h0000000000000100;
assign   tb_i_aad[926]                        =   tb_i_aad[925];
assign   tb_i_rf_static_plaintext_length[926] =   64'h0000000000000280;
assign   tb_i_plaintext[926]                  =   tb_i_plaintext[925];
assign   tb_o_valid[926]                      =   1'b0;
assign   tb_o_sop[926]                        =   1'b0;
assign   tb_o_ciphertext[926]                 =   tb_o_ciphertext[925];
assign   tb_o_tag_ready[926]                  =   1'b0;
assign   tb_o_tag[926]                        =   tb_o_tag[925];

// CLK no. 927/1240
// *************************************************
assign   tb_i_valid[927]                      =   1'b0;
assign   tb_i_reset[927]                      =   1'b0;
assign   tb_i_sop[927]                        =   1'b0;
assign   tb_i_key_update[927]                 =   1'b0;
assign   tb_i_key[927]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[927]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[927]               =   1'b0;
assign   tb_i_rf_static_encrypt[927]          =   1'b1;
assign   tb_i_clear_fault_flags[927]          =   1'b0;
assign   tb_i_rf_static_aad_length[927]       =   64'h0000000000000100;
assign   tb_i_aad[927]                        =   tb_i_aad[926];
assign   tb_i_rf_static_plaintext_length[927] =   64'h0000000000000280;
assign   tb_i_plaintext[927]                  =   tb_i_plaintext[926];
assign   tb_o_valid[927]                      =   1'b0;
assign   tb_o_sop[927]                        =   1'b0;
assign   tb_o_ciphertext[927]                 =   tb_o_ciphertext[926];
assign   tb_o_tag_ready[927]                  =   1'b0;
assign   tb_o_tag[927]                        =   tb_o_tag[926];

// CLK no. 928/1240
// *************************************************
assign   tb_i_valid[928]                      =   1'b0;
assign   tb_i_reset[928]                      =   1'b0;
assign   tb_i_sop[928]                        =   1'b0;
assign   tb_i_key_update[928]                 =   1'b0;
assign   tb_i_key[928]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[928]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[928]               =   1'b0;
assign   tb_i_rf_static_encrypt[928]          =   1'b1;
assign   tb_i_clear_fault_flags[928]          =   1'b0;
assign   tb_i_rf_static_aad_length[928]       =   64'h0000000000000100;
assign   tb_i_aad[928]                        =   tb_i_aad[927];
assign   tb_i_rf_static_plaintext_length[928] =   64'h0000000000000280;
assign   tb_i_plaintext[928]                  =   tb_i_plaintext[927];
assign   tb_o_valid[928]                      =   1'b0;
assign   tb_o_sop[928]                        =   1'b0;
assign   tb_o_ciphertext[928]                 =   tb_o_ciphertext[927];
assign   tb_o_tag_ready[928]                  =   1'b0;
assign   tb_o_tag[928]                        =   tb_o_tag[927];

// CLK no. 929/1240
// *************************************************
assign   tb_i_valid[929]                      =   1'b0;
assign   tb_i_reset[929]                      =   1'b0;
assign   tb_i_sop[929]                        =   1'b0;
assign   tb_i_key_update[929]                 =   1'b0;
assign   tb_i_key[929]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[929]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[929]               =   1'b0;
assign   tb_i_rf_static_encrypt[929]          =   1'b1;
assign   tb_i_clear_fault_flags[929]          =   1'b0;
assign   tb_i_rf_static_aad_length[929]       =   64'h0000000000000100;
assign   tb_i_aad[929]                        =   tb_i_aad[928];
assign   tb_i_rf_static_plaintext_length[929] =   64'h0000000000000280;
assign   tb_i_plaintext[929]                  =   tb_i_plaintext[928];
assign   tb_o_valid[929]                      =   1'b0;
assign   tb_o_sop[929]                        =   1'b0;
assign   tb_o_ciphertext[929]                 =   tb_o_ciphertext[928];
assign   tb_o_tag_ready[929]                  =   1'b0;
assign   tb_o_tag[929]                        =   tb_o_tag[928];

// CLK no. 930/1240
// *************************************************
assign   tb_i_valid[930]                      =   1'b0;
assign   tb_i_reset[930]                      =   1'b0;
assign   tb_i_sop[930]                        =   1'b0;
assign   tb_i_key_update[930]                 =   1'b0;
assign   tb_i_key[930]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[930]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[930]               =   1'b0;
assign   tb_i_rf_static_encrypt[930]          =   1'b1;
assign   tb_i_clear_fault_flags[930]          =   1'b0;
assign   tb_i_rf_static_aad_length[930]       =   64'h0000000000000100;
assign   tb_i_aad[930]                        =   tb_i_aad[929];
assign   tb_i_rf_static_plaintext_length[930] =   64'h0000000000000280;
assign   tb_i_plaintext[930]                  =   tb_i_plaintext[929];
assign   tb_o_valid[930]                      =   1'b0;
assign   tb_o_sop[930]                        =   1'b0;
assign   tb_o_ciphertext[930]                 =   tb_o_ciphertext[929];
assign   tb_o_tag_ready[930]                  =   1'b0;
assign   tb_o_tag[930]                        =   tb_o_tag[929];

// CLK no. 931/1240
// *************************************************
assign   tb_i_valid[931]                      =   1'b0;
assign   tb_i_reset[931]                      =   1'b0;
assign   tb_i_sop[931]                        =   1'b0;
assign   tb_i_key_update[931]                 =   1'b0;
assign   tb_i_key[931]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[931]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[931]               =   1'b0;
assign   tb_i_rf_static_encrypt[931]          =   1'b1;
assign   tb_i_clear_fault_flags[931]          =   1'b0;
assign   tb_i_rf_static_aad_length[931]       =   64'h0000000000000100;
assign   tb_i_aad[931]                        =   tb_i_aad[930];
assign   tb_i_rf_static_plaintext_length[931] =   64'h0000000000000280;
assign   tb_i_plaintext[931]                  =   tb_i_plaintext[930];
assign   tb_o_valid[931]                      =   1'b0;
assign   tb_o_sop[931]                        =   1'b0;
assign   tb_o_ciphertext[931]                 =   tb_o_ciphertext[930];
assign   tb_o_tag_ready[931]                  =   1'b0;
assign   tb_o_tag[931]                        =   tb_o_tag[930];

// CLK no. 932/1240
// *************************************************
assign   tb_i_valid[932]                      =   1'b0;
assign   tb_i_reset[932]                      =   1'b0;
assign   tb_i_sop[932]                        =   1'b0;
assign   tb_i_key_update[932]                 =   1'b0;
assign   tb_i_key[932]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[932]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[932]               =   1'b0;
assign   tb_i_rf_static_encrypt[932]          =   1'b1;
assign   tb_i_clear_fault_flags[932]          =   1'b0;
assign   tb_i_rf_static_aad_length[932]       =   64'h0000000000000100;
assign   tb_i_aad[932]                        =   tb_i_aad[931];
assign   tb_i_rf_static_plaintext_length[932] =   64'h0000000000000280;
assign   tb_i_plaintext[932]                  =   tb_i_plaintext[931];
assign   tb_o_valid[932]                      =   1'b1;
assign   tb_o_sop[932]                        =   1'b1;
assign   tb_o_ciphertext[932]                 =   256'hf179b589d25d0566361b3a4e5330e9a74ad29385b35fa11e169f3559875914f6;
assign   tb_o_tag_ready[932]                  =   1'b0;
assign   tb_o_tag[932]                        =   tb_o_tag[931];

// CLK no. 933/1240
// *************************************************
assign   tb_i_valid[933]                      =   1'b0;
assign   tb_i_reset[933]                      =   1'b0;
assign   tb_i_sop[933]                        =   1'b0;
assign   tb_i_key_update[933]                 =   1'b0;
assign   tb_i_key[933]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[933]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[933]               =   1'b0;
assign   tb_i_rf_static_encrypt[933]          =   1'b1;
assign   tb_i_clear_fault_flags[933]          =   1'b0;
assign   tb_i_rf_static_aad_length[933]       =   64'h0000000000000100;
assign   tb_i_aad[933]                        =   tb_i_aad[932];
assign   tb_i_rf_static_plaintext_length[933] =   64'h0000000000000280;
assign   tb_i_plaintext[933]                  =   tb_i_plaintext[932];
assign   tb_o_valid[933]                      =   1'b1;
assign   tb_o_sop[933]                        =   1'b0;
assign   tb_o_ciphertext[933]                 =   256'hca2a05cc6a620ee66c46a5b9a204667004aef481a23397ea2d6518219ea6c026;
assign   tb_o_tag_ready[933]                  =   1'b0;
assign   tb_o_tag[933]                        =   tb_o_tag[932];

// CLK no. 934/1240
// *************************************************
assign   tb_i_valid[934]                      =   1'b0;
assign   tb_i_reset[934]                      =   1'b0;
assign   tb_i_sop[934]                        =   1'b0;
assign   tb_i_key_update[934]                 =   1'b0;
assign   tb_i_key[934]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[934]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[934]               =   1'b0;
assign   tb_i_rf_static_encrypt[934]          =   1'b1;
assign   tb_i_clear_fault_flags[934]          =   1'b0;
assign   tb_i_rf_static_aad_length[934]       =   64'h0000000000000100;
assign   tb_i_aad[934]                        =   tb_i_aad[933];
assign   tb_i_rf_static_plaintext_length[934] =   64'h0000000000000280;
assign   tb_i_plaintext[934]                  =   tb_i_plaintext[933];
assign   tb_o_valid[934]                      =   1'b1;
assign   tb_o_sop[934]                        =   1'b0;
assign   tb_o_ciphertext[934]                 =   256'h6546af4795a7da30b4fd99f83e42eae8;
assign   tb_o_tag_ready[934]                  =   1'b0;
assign   tb_o_tag[934]                        =   tb_o_tag[933];

// CLK no. 935/1240
// *************************************************
assign   tb_i_valid[935]                      =   1'b0;
assign   tb_i_reset[935]                      =   1'b0;
assign   tb_i_sop[935]                        =   1'b0;
assign   tb_i_key_update[935]                 =   1'b0;
assign   tb_i_key[935]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[935]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[935]               =   1'b0;
assign   tb_i_rf_static_encrypt[935]          =   1'b1;
assign   tb_i_clear_fault_flags[935]          =   1'b0;
assign   tb_i_rf_static_aad_length[935]       =   64'h0000000000000100;
assign   tb_i_aad[935]                        =   tb_i_aad[934];
assign   tb_i_rf_static_plaintext_length[935] =   64'h0000000000000280;
assign   tb_i_plaintext[935]                  =   tb_i_plaintext[934];
assign   tb_o_valid[935]                      =   1'b0;
assign   tb_o_sop[935]                        =   1'b0;
assign   tb_o_ciphertext[935]                 =   tb_o_ciphertext[934];
assign   tb_o_tag_ready[935]                  =   1'b0;
assign   tb_o_tag[935]                        =   tb_o_tag[934];

// CLK no. 936/1240
// *************************************************
assign   tb_i_valid[936]                      =   1'b0;
assign   tb_i_reset[936]                      =   1'b0;
assign   tb_i_sop[936]                        =   1'b0;
assign   tb_i_key_update[936]                 =   1'b0;
assign   tb_i_key[936]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[936]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[936]               =   1'b0;
assign   tb_i_rf_static_encrypt[936]          =   1'b1;
assign   tb_i_clear_fault_flags[936]          =   1'b0;
assign   tb_i_rf_static_aad_length[936]       =   64'h0000000000000100;
assign   tb_i_aad[936]                        =   tb_i_aad[935];
assign   tb_i_rf_static_plaintext_length[936] =   64'h0000000000000280;
assign   tb_i_plaintext[936]                  =   tb_i_plaintext[935];
assign   tb_o_valid[936]                      =   1'b0;
assign   tb_o_sop[936]                        =   1'b0;
assign   tb_o_ciphertext[936]                 =   tb_o_ciphertext[935];
assign   tb_o_tag_ready[936]                  =   1'b0;
assign   tb_o_tag[936]                        =   tb_o_tag[935];

// CLK no. 937/1240
// *************************************************
assign   tb_i_valid[937]                      =   1'b0;
assign   tb_i_reset[937]                      =   1'b0;
assign   tb_i_sop[937]                        =   1'b0;
assign   tb_i_key_update[937]                 =   1'b0;
assign   tb_i_key[937]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[937]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[937]               =   1'b0;
assign   tb_i_rf_static_encrypt[937]          =   1'b1;
assign   tb_i_clear_fault_flags[937]          =   1'b0;
assign   tb_i_rf_static_aad_length[937]       =   64'h0000000000000100;
assign   tb_i_aad[937]                        =   tb_i_aad[936];
assign   tb_i_rf_static_plaintext_length[937] =   64'h0000000000000280;
assign   tb_i_plaintext[937]                  =   tb_i_plaintext[936];
assign   tb_o_valid[937]                      =   1'b0;
assign   tb_o_sop[937]                        =   1'b0;
assign   tb_o_ciphertext[937]                 =   tb_o_ciphertext[936];
assign   tb_o_tag_ready[937]                  =   1'b0;
assign   tb_o_tag[937]                        =   tb_o_tag[936];

// CLK no. 938/1240
// *************************************************
assign   tb_i_valid[938]                      =   1'b0;
assign   tb_i_reset[938]                      =   1'b0;
assign   tb_i_sop[938]                        =   1'b0;
assign   tb_i_key_update[938]                 =   1'b0;
assign   tb_i_key[938]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[938]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[938]               =   1'b0;
assign   tb_i_rf_static_encrypt[938]          =   1'b1;
assign   tb_i_clear_fault_flags[938]          =   1'b0;
assign   tb_i_rf_static_aad_length[938]       =   64'h0000000000000100;
assign   tb_i_aad[938]                        =   tb_i_aad[937];
assign   tb_i_rf_static_plaintext_length[938] =   64'h0000000000000280;
assign   tb_i_plaintext[938]                  =   tb_i_plaintext[937];
assign   tb_o_valid[938]                      =   1'b0;
assign   tb_o_sop[938]                        =   1'b0;
assign   tb_o_ciphertext[938]                 =   tb_o_ciphertext[937];
assign   tb_o_tag_ready[938]                  =   1'b0;
assign   tb_o_tag[938]                        =   tb_o_tag[937];

// CLK no. 939/1240
// *************************************************
assign   tb_i_valid[939]                      =   1'b0;
assign   tb_i_reset[939]                      =   1'b0;
assign   tb_i_sop[939]                        =   1'b0;
assign   tb_i_key_update[939]                 =   1'b0;
assign   tb_i_key[939]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[939]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[939]               =   1'b0;
assign   tb_i_rf_static_encrypt[939]          =   1'b1;
assign   tb_i_clear_fault_flags[939]          =   1'b0;
assign   tb_i_rf_static_aad_length[939]       =   64'h0000000000000100;
assign   tb_i_aad[939]                        =   tb_i_aad[938];
assign   tb_i_rf_static_plaintext_length[939] =   64'h0000000000000280;
assign   tb_i_plaintext[939]                  =   tb_i_plaintext[938];
assign   tb_o_valid[939]                      =   1'b0;
assign   tb_o_sop[939]                        =   1'b0;
assign   tb_o_ciphertext[939]                 =   tb_o_ciphertext[938];
assign   tb_o_tag_ready[939]                  =   1'b0;
assign   tb_o_tag[939]                        =   tb_o_tag[938];

// CLK no. 940/1240
// *************************************************
assign   tb_i_valid[940]                      =   1'b0;
assign   tb_i_reset[940]                      =   1'b0;
assign   tb_i_sop[940]                        =   1'b0;
assign   tb_i_key_update[940]                 =   1'b0;
assign   tb_i_key[940]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[940]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[940]               =   1'b0;
assign   tb_i_rf_static_encrypt[940]          =   1'b1;
assign   tb_i_clear_fault_flags[940]          =   1'b0;
assign   tb_i_rf_static_aad_length[940]       =   64'h0000000000000100;
assign   tb_i_aad[940]                        =   tb_i_aad[939];
assign   tb_i_rf_static_plaintext_length[940] =   64'h0000000000000280;
assign   tb_i_plaintext[940]                  =   tb_i_plaintext[939];
assign   tb_o_valid[940]                      =   1'b0;
assign   tb_o_sop[940]                        =   1'b0;
assign   tb_o_ciphertext[940]                 =   tb_o_ciphertext[939];
assign   tb_o_tag_ready[940]                  =   1'b0;
assign   tb_o_tag[940]                        =   tb_o_tag[939];

// CLK no. 941/1240
// *************************************************
assign   tb_i_valid[941]                      =   1'b0;
assign   tb_i_reset[941]                      =   1'b0;
assign   tb_i_sop[941]                        =   1'b0;
assign   tb_i_key_update[941]                 =   1'b0;
assign   tb_i_key[941]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[941]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[941]               =   1'b0;
assign   tb_i_rf_static_encrypt[941]          =   1'b1;
assign   tb_i_clear_fault_flags[941]          =   1'b0;
assign   tb_i_rf_static_aad_length[941]       =   64'h0000000000000100;
assign   tb_i_aad[941]                        =   tb_i_aad[940];
assign   tb_i_rf_static_plaintext_length[941] =   64'h0000000000000280;
assign   tb_i_plaintext[941]                  =   tb_i_plaintext[940];
assign   tb_o_valid[941]                      =   1'b0;
assign   tb_o_sop[941]                        =   1'b0;
assign   tb_o_ciphertext[941]                 =   tb_o_ciphertext[940];
assign   tb_o_tag_ready[941]                  =   1'b0;
assign   tb_o_tag[941]                        =   tb_o_tag[940];

// CLK no. 942/1240
// *************************************************
assign   tb_i_valid[942]                      =   1'b0;
assign   tb_i_reset[942]                      =   1'b0;
assign   tb_i_sop[942]                        =   1'b0;
assign   tb_i_key_update[942]                 =   1'b0;
assign   tb_i_key[942]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[942]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[942]               =   1'b0;
assign   tb_i_rf_static_encrypt[942]          =   1'b1;
assign   tb_i_clear_fault_flags[942]          =   1'b0;
assign   tb_i_rf_static_aad_length[942]       =   64'h0000000000000100;
assign   tb_i_aad[942]                        =   tb_i_aad[941];
assign   tb_i_rf_static_plaintext_length[942] =   64'h0000000000000280;
assign   tb_i_plaintext[942]                  =   tb_i_plaintext[941];
assign   tb_o_valid[942]                      =   1'b0;
assign   tb_o_sop[942]                        =   1'b0;
assign   tb_o_ciphertext[942]                 =   tb_o_ciphertext[941];
assign   tb_o_tag_ready[942]                  =   1'b1;
assign   tb_o_tag[942]                        =   128'hb2b203b38875e696a033633f6d58ba9c;

// CLK no. 943/1240
// *************************************************
assign   tb_i_valid[943]                      =   1'b0;
assign   tb_i_reset[943]                      =   1'b0;
assign   tb_i_sop[943]                        =   1'b0;
assign   tb_i_key_update[943]                 =   1'b0;
assign   tb_i_key[943]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[943]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[943]               =   1'b0;
assign   tb_i_rf_static_encrypt[943]          =   1'b1;
assign   tb_i_clear_fault_flags[943]          =   1'b0;
assign   tb_i_rf_static_aad_length[943]       =   64'h0000000000000100;
assign   tb_i_aad[943]                        =   tb_i_aad[942];
assign   tb_i_rf_static_plaintext_length[943] =   64'h0000000000000280;
assign   tb_i_plaintext[943]                  =   tb_i_plaintext[942];
assign   tb_o_valid[943]                      =   1'b0;
assign   tb_o_sop[943]                        =   1'b0;
assign   tb_o_ciphertext[943]                 =   tb_o_ciphertext[942];
assign   tb_o_tag_ready[943]                  =   1'b0;
assign   tb_o_tag[943]                        =   tb_o_tag[942];

// CLK no. 944/1240
// *************************************************
assign   tb_i_valid[944]                      =   1'b0;
assign   tb_i_reset[944]                      =   1'b0;
assign   tb_i_sop[944]                        =   1'b0;
assign   tb_i_key_update[944]                 =   1'b0;
assign   tb_i_key[944]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[944]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[944]               =   1'b0;
assign   tb_i_rf_static_encrypt[944]          =   1'b1;
assign   tb_i_clear_fault_flags[944]          =   1'b0;
assign   tb_i_rf_static_aad_length[944]       =   64'h0000000000000100;
assign   tb_i_aad[944]                        =   tb_i_aad[943];
assign   tb_i_rf_static_plaintext_length[944] =   64'h0000000000000280;
assign   tb_i_plaintext[944]                  =   tb_i_plaintext[943];
assign   tb_o_valid[944]                      =   1'b0;
assign   tb_o_sop[944]                        =   1'b0;
assign   tb_o_ciphertext[944]                 =   tb_o_ciphertext[943];
assign   tb_o_tag_ready[944]                  =   1'b0;
assign   tb_o_tag[944]                        =   tb_o_tag[943];

// CLK no. 945/1240
// *************************************************
assign   tb_i_valid[945]                      =   1'b0;
assign   tb_i_reset[945]                      =   1'b0;
assign   tb_i_sop[945]                        =   1'b1;
assign   tb_i_key_update[945]                 =   1'b0;
assign   tb_i_key[945]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[945]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[945]               =   1'b0;
assign   tb_i_rf_static_encrypt[945]          =   1'b1;
assign   tb_i_clear_fault_flags[945]          =   1'b0;
assign   tb_i_rf_static_aad_length[945]       =   64'h0000000000000100;
assign   tb_i_aad[945]                        =   tb_i_aad[944];
assign   tb_i_rf_static_plaintext_length[945] =   64'h0000000000000280;
assign   tb_i_plaintext[945]                  =   tb_i_plaintext[944];
assign   tb_o_valid[945]                      =   1'b0;
assign   tb_o_sop[945]                        =   1'b0;
assign   tb_o_ciphertext[945]                 =   tb_o_ciphertext[944];
assign   tb_o_tag_ready[945]                  =   1'b0;
assign   tb_o_tag[945]                        =   tb_o_tag[944];

// CLK no. 946/1240
// *************************************************
assign   tb_i_valid[946]                      =   1'b1;
assign   tb_i_reset[946]                      =   1'b0;
assign   tb_i_sop[946]                        =   1'b0;
assign   tb_i_key_update[946]                 =   1'b0;
assign   tb_i_key[946]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[946]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[946]               =   1'b0;
assign   tb_i_rf_static_encrypt[946]          =   1'b1;
assign   tb_i_clear_fault_flags[946]          =   1'b0;
assign   tb_i_rf_static_aad_length[946]       =   64'h0000000000000100;
assign   tb_i_aad[946]                        =   256'h81deddab3b9a4e2880fe7000f2b3f1abb1c5d6c14fa8457b48b55dda3e83ff1c;
assign   tb_i_rf_static_plaintext_length[946] =   64'h0000000000000280;
assign   tb_i_plaintext[946]                  =   tb_i_plaintext[945];
assign   tb_o_valid[946]                      =   1'b0;
assign   tb_o_sop[946]                        =   1'b0;
assign   tb_o_ciphertext[946]                 =   tb_o_ciphertext[945];
assign   tb_o_tag_ready[946]                  =   1'b0;
assign   tb_o_tag[946]                        =   tb_o_tag[945];

// CLK no. 947/1240
// *************************************************
assign   tb_i_valid[947]                      =   1'b1;
assign   tb_i_reset[947]                      =   1'b0;
assign   tb_i_sop[947]                        =   1'b0;
assign   tb_i_key_update[947]                 =   1'b0;
assign   tb_i_key[947]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[947]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[947]               =   1'b0;
assign   tb_i_rf_static_encrypt[947]          =   1'b1;
assign   tb_i_clear_fault_flags[947]          =   1'b0;
assign   tb_i_rf_static_aad_length[947]       =   64'h0000000000000100;
assign   tb_i_aad[947]                        =   tb_i_aad[946];
assign   tb_i_rf_static_plaintext_length[947] =   64'h0000000000000280;
assign   tb_i_plaintext[947]                  =   256'haa03596f1389f41191c80e18defdf31a90b32ff4fea5d381640b309a6423d4af;
assign   tb_o_valid[947]                      =   1'b0;
assign   tb_o_sop[947]                        =   1'b0;
assign   tb_o_ciphertext[947]                 =   tb_o_ciphertext[946];
assign   tb_o_tag_ready[947]                  =   1'b0;
assign   tb_o_tag[947]                        =   tb_o_tag[946];

// CLK no. 948/1240
// *************************************************
assign   tb_i_valid[948]                      =   1'b1;
assign   tb_i_reset[948]                      =   1'b0;
assign   tb_i_sop[948]                        =   1'b0;
assign   tb_i_key_update[948]                 =   1'b0;
assign   tb_i_key[948]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[948]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[948]               =   1'b0;
assign   tb_i_rf_static_encrypt[948]          =   1'b1;
assign   tb_i_clear_fault_flags[948]          =   1'b0;
assign   tb_i_rf_static_aad_length[948]       =   64'h0000000000000100;
assign   tb_i_aad[948]                        =   tb_i_aad[947];
assign   tb_i_rf_static_plaintext_length[948] =   64'h0000000000000280;
assign   tb_i_plaintext[948]                  =   256'hecd6a0c4bfc06ddeed5088a1484fcc797162676d9562d6a5e1761ac86cc67da2;
assign   tb_o_valid[948]                      =   1'b0;
assign   tb_o_sop[948]                        =   1'b0;
assign   tb_o_ciphertext[948]                 =   tb_o_ciphertext[947];
assign   tb_o_tag_ready[948]                  =   1'b0;
assign   tb_o_tag[948]                        =   tb_o_tag[947];

// CLK no. 949/1240
// *************************************************
assign   tb_i_valid[949]                      =   1'b1;
assign   tb_i_reset[949]                      =   1'b0;
assign   tb_i_sop[949]                        =   1'b0;
assign   tb_i_key_update[949]                 =   1'b0;
assign   tb_i_key[949]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[949]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[949]               =   1'b0;
assign   tb_i_rf_static_encrypt[949]          =   1'b1;
assign   tb_i_clear_fault_flags[949]          =   1'b0;
assign   tb_i_rf_static_aad_length[949]       =   64'h0000000000000100;
assign   tb_i_aad[949]                        =   tb_i_aad[948];
assign   tb_i_rf_static_plaintext_length[949] =   64'h0000000000000280;
assign   tb_i_plaintext[949]                  =   256'h494b75040e115f71b2884ec4f0063844;
assign   tb_o_valid[949]                      =   1'b0;
assign   tb_o_sop[949]                        =   1'b0;
assign   tb_o_ciphertext[949]                 =   tb_o_ciphertext[948];
assign   tb_o_tag_ready[949]                  =   1'b0;
assign   tb_o_tag[949]                        =   tb_o_tag[948];

// CLK no. 950/1240
// *************************************************
assign   tb_i_valid[950]                      =   1'b0;
assign   tb_i_reset[950]                      =   1'b0;
assign   tb_i_sop[950]                        =   1'b0;
assign   tb_i_key_update[950]                 =   1'b0;
assign   tb_i_key[950]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[950]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[950]               =   1'b0;
assign   tb_i_rf_static_encrypt[950]          =   1'b1;
assign   tb_i_clear_fault_flags[950]          =   1'b0;
assign   tb_i_rf_static_aad_length[950]       =   64'h0000000000000100;
assign   tb_i_aad[950]                        =   tb_i_aad[949];
assign   tb_i_rf_static_plaintext_length[950] =   64'h0000000000000280;
assign   tb_i_plaintext[950]                  =   tb_i_plaintext[949];
assign   tb_o_valid[950]                      =   1'b0;
assign   tb_o_sop[950]                        =   1'b0;
assign   tb_o_ciphertext[950]                 =   tb_o_ciphertext[949];
assign   tb_o_tag_ready[950]                  =   1'b0;
assign   tb_o_tag[950]                        =   tb_o_tag[949];

// CLK no. 951/1240
// *************************************************
assign   tb_i_valid[951]                      =   1'b0;
assign   tb_i_reset[951]                      =   1'b0;
assign   tb_i_sop[951]                        =   1'b0;
assign   tb_i_key_update[951]                 =   1'b0;
assign   tb_i_key[951]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[951]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[951]               =   1'b0;
assign   tb_i_rf_static_encrypt[951]          =   1'b1;
assign   tb_i_clear_fault_flags[951]          =   1'b0;
assign   tb_i_rf_static_aad_length[951]       =   64'h0000000000000100;
assign   tb_i_aad[951]                        =   tb_i_aad[950];
assign   tb_i_rf_static_plaintext_length[951] =   64'h0000000000000280;
assign   tb_i_plaintext[951]                  =   tb_i_plaintext[950];
assign   tb_o_valid[951]                      =   1'b0;
assign   tb_o_sop[951]                        =   1'b0;
assign   tb_o_ciphertext[951]                 =   tb_o_ciphertext[950];
assign   tb_o_tag_ready[951]                  =   1'b0;
assign   tb_o_tag[951]                        =   tb_o_tag[950];

// CLK no. 952/1240
// *************************************************
assign   tb_i_valid[952]                      =   1'b0;
assign   tb_i_reset[952]                      =   1'b0;
assign   tb_i_sop[952]                        =   1'b0;
assign   tb_i_key_update[952]                 =   1'b0;
assign   tb_i_key[952]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[952]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[952]               =   1'b0;
assign   tb_i_rf_static_encrypt[952]          =   1'b1;
assign   tb_i_clear_fault_flags[952]          =   1'b0;
assign   tb_i_rf_static_aad_length[952]       =   64'h0000000000000100;
assign   tb_i_aad[952]                        =   tb_i_aad[951];
assign   tb_i_rf_static_plaintext_length[952] =   64'h0000000000000280;
assign   tb_i_plaintext[952]                  =   tb_i_plaintext[951];
assign   tb_o_valid[952]                      =   1'b0;
assign   tb_o_sop[952]                        =   1'b0;
assign   tb_o_ciphertext[952]                 =   tb_o_ciphertext[951];
assign   tb_o_tag_ready[952]                  =   1'b0;
assign   tb_o_tag[952]                        =   tb_o_tag[951];

// CLK no. 953/1240
// *************************************************
assign   tb_i_valid[953]                      =   1'b0;
assign   tb_i_reset[953]                      =   1'b0;
assign   tb_i_sop[953]                        =   1'b0;
assign   tb_i_key_update[953]                 =   1'b0;
assign   tb_i_key[953]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[953]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[953]               =   1'b0;
assign   tb_i_rf_static_encrypt[953]          =   1'b1;
assign   tb_i_clear_fault_flags[953]          =   1'b0;
assign   tb_i_rf_static_aad_length[953]       =   64'h0000000000000100;
assign   tb_i_aad[953]                        =   tb_i_aad[952];
assign   tb_i_rf_static_plaintext_length[953] =   64'h0000000000000280;
assign   tb_i_plaintext[953]                  =   tb_i_plaintext[952];
assign   tb_o_valid[953]                      =   1'b0;
assign   tb_o_sop[953]                        =   1'b0;
assign   tb_o_ciphertext[953]                 =   tb_o_ciphertext[952];
assign   tb_o_tag_ready[953]                  =   1'b0;
assign   tb_o_tag[953]                        =   tb_o_tag[952];

// CLK no. 954/1240
// *************************************************
assign   tb_i_valid[954]                      =   1'b0;
assign   tb_i_reset[954]                      =   1'b0;
assign   tb_i_sop[954]                        =   1'b0;
assign   tb_i_key_update[954]                 =   1'b0;
assign   tb_i_key[954]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[954]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[954]               =   1'b0;
assign   tb_i_rf_static_encrypt[954]          =   1'b1;
assign   tb_i_clear_fault_flags[954]          =   1'b0;
assign   tb_i_rf_static_aad_length[954]       =   64'h0000000000000100;
assign   tb_i_aad[954]                        =   tb_i_aad[953];
assign   tb_i_rf_static_plaintext_length[954] =   64'h0000000000000280;
assign   tb_i_plaintext[954]                  =   tb_i_plaintext[953];
assign   tb_o_valid[954]                      =   1'b0;
assign   tb_o_sop[954]                        =   1'b0;
assign   tb_o_ciphertext[954]                 =   tb_o_ciphertext[953];
assign   tb_o_tag_ready[954]                  =   1'b0;
assign   tb_o_tag[954]                        =   tb_o_tag[953];

// CLK no. 955/1240
// *************************************************
assign   tb_i_valid[955]                      =   1'b0;
assign   tb_i_reset[955]                      =   1'b0;
assign   tb_i_sop[955]                        =   1'b0;
assign   tb_i_key_update[955]                 =   1'b0;
assign   tb_i_key[955]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[955]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[955]               =   1'b0;
assign   tb_i_rf_static_encrypt[955]          =   1'b1;
assign   tb_i_clear_fault_flags[955]          =   1'b0;
assign   tb_i_rf_static_aad_length[955]       =   64'h0000000000000100;
assign   tb_i_aad[955]                        =   tb_i_aad[954];
assign   tb_i_rf_static_plaintext_length[955] =   64'h0000000000000280;
assign   tb_i_plaintext[955]                  =   tb_i_plaintext[954];
assign   tb_o_valid[955]                      =   1'b0;
assign   tb_o_sop[955]                        =   1'b0;
assign   tb_o_ciphertext[955]                 =   tb_o_ciphertext[954];
assign   tb_o_tag_ready[955]                  =   1'b0;
assign   tb_o_tag[955]                        =   tb_o_tag[954];

// CLK no. 956/1240
// *************************************************
assign   tb_i_valid[956]                      =   1'b0;
assign   tb_i_reset[956]                      =   1'b0;
assign   tb_i_sop[956]                        =   1'b0;
assign   tb_i_key_update[956]                 =   1'b0;
assign   tb_i_key[956]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[956]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[956]               =   1'b0;
assign   tb_i_rf_static_encrypt[956]          =   1'b1;
assign   tb_i_clear_fault_flags[956]          =   1'b0;
assign   tb_i_rf_static_aad_length[956]       =   64'h0000000000000100;
assign   tb_i_aad[956]                        =   tb_i_aad[955];
assign   tb_i_rf_static_plaintext_length[956] =   64'h0000000000000280;
assign   tb_i_plaintext[956]                  =   tb_i_plaintext[955];
assign   tb_o_valid[956]                      =   1'b0;
assign   tb_o_sop[956]                        =   1'b0;
assign   tb_o_ciphertext[956]                 =   tb_o_ciphertext[955];
assign   tb_o_tag_ready[956]                  =   1'b0;
assign   tb_o_tag[956]                        =   tb_o_tag[955];

// CLK no. 957/1240
// *************************************************
assign   tb_i_valid[957]                      =   1'b0;
assign   tb_i_reset[957]                      =   1'b0;
assign   tb_i_sop[957]                        =   1'b0;
assign   tb_i_key_update[957]                 =   1'b0;
assign   tb_i_key[957]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[957]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[957]               =   1'b0;
assign   tb_i_rf_static_encrypt[957]          =   1'b1;
assign   tb_i_clear_fault_flags[957]          =   1'b0;
assign   tb_i_rf_static_aad_length[957]       =   64'h0000000000000100;
assign   tb_i_aad[957]                        =   tb_i_aad[956];
assign   tb_i_rf_static_plaintext_length[957] =   64'h0000000000000280;
assign   tb_i_plaintext[957]                  =   tb_i_plaintext[956];
assign   tb_o_valid[957]                      =   1'b0;
assign   tb_o_sop[957]                        =   1'b0;
assign   tb_o_ciphertext[957]                 =   tb_o_ciphertext[956];
assign   tb_o_tag_ready[957]                  =   1'b0;
assign   tb_o_tag[957]                        =   tb_o_tag[956];

// CLK no. 958/1240
// *************************************************
assign   tb_i_valid[958]                      =   1'b0;
assign   tb_i_reset[958]                      =   1'b0;
assign   tb_i_sop[958]                        =   1'b0;
assign   tb_i_key_update[958]                 =   1'b0;
assign   tb_i_key[958]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[958]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[958]               =   1'b0;
assign   tb_i_rf_static_encrypt[958]          =   1'b1;
assign   tb_i_clear_fault_flags[958]          =   1'b0;
assign   tb_i_rf_static_aad_length[958]       =   64'h0000000000000100;
assign   tb_i_aad[958]                        =   tb_i_aad[957];
assign   tb_i_rf_static_plaintext_length[958] =   64'h0000000000000280;
assign   tb_i_plaintext[958]                  =   tb_i_plaintext[957];
assign   tb_o_valid[958]                      =   1'b0;
assign   tb_o_sop[958]                        =   1'b0;
assign   tb_o_ciphertext[958]                 =   tb_o_ciphertext[957];
assign   tb_o_tag_ready[958]                  =   1'b0;
assign   tb_o_tag[958]                        =   tb_o_tag[957];

// CLK no. 959/1240
// *************************************************
assign   tb_i_valid[959]                      =   1'b0;
assign   tb_i_reset[959]                      =   1'b0;
assign   tb_i_sop[959]                        =   1'b0;
assign   tb_i_key_update[959]                 =   1'b0;
assign   tb_i_key[959]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[959]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[959]               =   1'b0;
assign   tb_i_rf_static_encrypt[959]          =   1'b1;
assign   tb_i_clear_fault_flags[959]          =   1'b0;
assign   tb_i_rf_static_aad_length[959]       =   64'h0000000000000100;
assign   tb_i_aad[959]                        =   tb_i_aad[958];
assign   tb_i_rf_static_plaintext_length[959] =   64'h0000000000000280;
assign   tb_i_plaintext[959]                  =   tb_i_plaintext[958];
assign   tb_o_valid[959]                      =   1'b0;
assign   tb_o_sop[959]                        =   1'b0;
assign   tb_o_ciphertext[959]                 =   tb_o_ciphertext[958];
assign   tb_o_tag_ready[959]                  =   1'b0;
assign   tb_o_tag[959]                        =   tb_o_tag[958];

// CLK no. 960/1240
// *************************************************
assign   tb_i_valid[960]                      =   1'b0;
assign   tb_i_reset[960]                      =   1'b0;
assign   tb_i_sop[960]                        =   1'b0;
assign   tb_i_key_update[960]                 =   1'b0;
assign   tb_i_key[960]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[960]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[960]               =   1'b0;
assign   tb_i_rf_static_encrypt[960]          =   1'b1;
assign   tb_i_clear_fault_flags[960]          =   1'b0;
assign   tb_i_rf_static_aad_length[960]       =   64'h0000000000000100;
assign   tb_i_aad[960]                        =   tb_i_aad[959];
assign   tb_i_rf_static_plaintext_length[960] =   64'h0000000000000280;
assign   tb_i_plaintext[960]                  =   tb_i_plaintext[959];
assign   tb_o_valid[960]                      =   1'b0;
assign   tb_o_sop[960]                        =   1'b0;
assign   tb_o_ciphertext[960]                 =   tb_o_ciphertext[959];
assign   tb_o_tag_ready[960]                  =   1'b0;
assign   tb_o_tag[960]                        =   tb_o_tag[959];

// CLK no. 961/1240
// *************************************************
assign   tb_i_valid[961]                      =   1'b0;
assign   tb_i_reset[961]                      =   1'b0;
assign   tb_i_sop[961]                        =   1'b0;
assign   tb_i_key_update[961]                 =   1'b0;
assign   tb_i_key[961]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[961]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[961]               =   1'b0;
assign   tb_i_rf_static_encrypt[961]          =   1'b1;
assign   tb_i_clear_fault_flags[961]          =   1'b0;
assign   tb_i_rf_static_aad_length[961]       =   64'h0000000000000100;
assign   tb_i_aad[961]                        =   tb_i_aad[960];
assign   tb_i_rf_static_plaintext_length[961] =   64'h0000000000000280;
assign   tb_i_plaintext[961]                  =   tb_i_plaintext[960];
assign   tb_o_valid[961]                      =   1'b0;
assign   tb_o_sop[961]                        =   1'b0;
assign   tb_o_ciphertext[961]                 =   tb_o_ciphertext[960];
assign   tb_o_tag_ready[961]                  =   1'b0;
assign   tb_o_tag[961]                        =   tb_o_tag[960];

// CLK no. 962/1240
// *************************************************
assign   tb_i_valid[962]                      =   1'b0;
assign   tb_i_reset[962]                      =   1'b0;
assign   tb_i_sop[962]                        =   1'b0;
assign   tb_i_key_update[962]                 =   1'b0;
assign   tb_i_key[962]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[962]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[962]               =   1'b0;
assign   tb_i_rf_static_encrypt[962]          =   1'b1;
assign   tb_i_clear_fault_flags[962]          =   1'b0;
assign   tb_i_rf_static_aad_length[962]       =   64'h0000000000000100;
assign   tb_i_aad[962]                        =   tb_i_aad[961];
assign   tb_i_rf_static_plaintext_length[962] =   64'h0000000000000280;
assign   tb_i_plaintext[962]                  =   tb_i_plaintext[961];
assign   tb_o_valid[962]                      =   1'b0;
assign   tb_o_sop[962]                        =   1'b0;
assign   tb_o_ciphertext[962]                 =   tb_o_ciphertext[961];
assign   tb_o_tag_ready[962]                  =   1'b0;
assign   tb_o_tag[962]                        =   tb_o_tag[961];

// CLK no. 963/1240
// *************************************************
assign   tb_i_valid[963]                      =   1'b0;
assign   tb_i_reset[963]                      =   1'b0;
assign   tb_i_sop[963]                        =   1'b0;
assign   tb_i_key_update[963]                 =   1'b0;
assign   tb_i_key[963]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[963]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[963]               =   1'b0;
assign   tb_i_rf_static_encrypt[963]          =   1'b1;
assign   tb_i_clear_fault_flags[963]          =   1'b0;
assign   tb_i_rf_static_aad_length[963]       =   64'h0000000000000100;
assign   tb_i_aad[963]                        =   tb_i_aad[962];
assign   tb_i_rf_static_plaintext_length[963] =   64'h0000000000000280;
assign   tb_i_plaintext[963]                  =   tb_i_plaintext[962];
assign   tb_o_valid[963]                      =   1'b0;
assign   tb_o_sop[963]                        =   1'b0;
assign   tb_o_ciphertext[963]                 =   tb_o_ciphertext[962];
assign   tb_o_tag_ready[963]                  =   1'b0;
assign   tb_o_tag[963]                        =   tb_o_tag[962];

// CLK no. 964/1240
// *************************************************
assign   tb_i_valid[964]                      =   1'b0;
assign   tb_i_reset[964]                      =   1'b0;
assign   tb_i_sop[964]                        =   1'b0;
assign   tb_i_key_update[964]                 =   1'b0;
assign   tb_i_key[964]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[964]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[964]               =   1'b0;
assign   tb_i_rf_static_encrypt[964]          =   1'b1;
assign   tb_i_clear_fault_flags[964]          =   1'b0;
assign   tb_i_rf_static_aad_length[964]       =   64'h0000000000000100;
assign   tb_i_aad[964]                        =   tb_i_aad[963];
assign   tb_i_rf_static_plaintext_length[964] =   64'h0000000000000280;
assign   tb_i_plaintext[964]                  =   tb_i_plaintext[963];
assign   tb_o_valid[964]                      =   1'b0;
assign   tb_o_sop[964]                        =   1'b0;
assign   tb_o_ciphertext[964]                 =   tb_o_ciphertext[963];
assign   tb_o_tag_ready[964]                  =   1'b0;
assign   tb_o_tag[964]                        =   tb_o_tag[963];

// CLK no. 965/1240
// *************************************************
assign   tb_i_valid[965]                      =   1'b0;
assign   tb_i_reset[965]                      =   1'b0;
assign   tb_i_sop[965]                        =   1'b0;
assign   tb_i_key_update[965]                 =   1'b0;
assign   tb_i_key[965]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[965]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[965]               =   1'b0;
assign   tb_i_rf_static_encrypt[965]          =   1'b1;
assign   tb_i_clear_fault_flags[965]          =   1'b0;
assign   tb_i_rf_static_aad_length[965]       =   64'h0000000000000100;
assign   tb_i_aad[965]                        =   tb_i_aad[964];
assign   tb_i_rf_static_plaintext_length[965] =   64'h0000000000000280;
assign   tb_i_plaintext[965]                  =   tb_i_plaintext[964];
assign   tb_o_valid[965]                      =   1'b0;
assign   tb_o_sop[965]                        =   1'b0;
assign   tb_o_ciphertext[965]                 =   tb_o_ciphertext[964];
assign   tb_o_tag_ready[965]                  =   1'b0;
assign   tb_o_tag[965]                        =   tb_o_tag[964];

// CLK no. 966/1240
// *************************************************
assign   tb_i_valid[966]                      =   1'b0;
assign   tb_i_reset[966]                      =   1'b0;
assign   tb_i_sop[966]                        =   1'b0;
assign   tb_i_key_update[966]                 =   1'b0;
assign   tb_i_key[966]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[966]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[966]               =   1'b0;
assign   tb_i_rf_static_encrypt[966]          =   1'b1;
assign   tb_i_clear_fault_flags[966]          =   1'b0;
assign   tb_i_rf_static_aad_length[966]       =   64'h0000000000000100;
assign   tb_i_aad[966]                        =   tb_i_aad[965];
assign   tb_i_rf_static_plaintext_length[966] =   64'h0000000000000280;
assign   tb_i_plaintext[966]                  =   tb_i_plaintext[965];
assign   tb_o_valid[966]                      =   1'b0;
assign   tb_o_sop[966]                        =   1'b0;
assign   tb_o_ciphertext[966]                 =   tb_o_ciphertext[965];
assign   tb_o_tag_ready[966]                  =   1'b0;
assign   tb_o_tag[966]                        =   tb_o_tag[965];

// CLK no. 967/1240
// *************************************************
assign   tb_i_valid[967]                      =   1'b0;
assign   tb_i_reset[967]                      =   1'b0;
assign   tb_i_sop[967]                        =   1'b0;
assign   tb_i_key_update[967]                 =   1'b0;
assign   tb_i_key[967]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[967]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[967]               =   1'b0;
assign   tb_i_rf_static_encrypt[967]          =   1'b1;
assign   tb_i_clear_fault_flags[967]          =   1'b0;
assign   tb_i_rf_static_aad_length[967]       =   64'h0000000000000100;
assign   tb_i_aad[967]                        =   tb_i_aad[966];
assign   tb_i_rf_static_plaintext_length[967] =   64'h0000000000000280;
assign   tb_i_plaintext[967]                  =   tb_i_plaintext[966];
assign   tb_o_valid[967]                      =   1'b0;
assign   tb_o_sop[967]                        =   1'b0;
assign   tb_o_ciphertext[967]                 =   tb_o_ciphertext[966];
assign   tb_o_tag_ready[967]                  =   1'b0;
assign   tb_o_tag[967]                        =   tb_o_tag[966];

// CLK no. 968/1240
// *************************************************
assign   tb_i_valid[968]                      =   1'b0;
assign   tb_i_reset[968]                      =   1'b0;
assign   tb_i_sop[968]                        =   1'b0;
assign   tb_i_key_update[968]                 =   1'b0;
assign   tb_i_key[968]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[968]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[968]               =   1'b0;
assign   tb_i_rf_static_encrypt[968]          =   1'b1;
assign   tb_i_clear_fault_flags[968]          =   1'b0;
assign   tb_i_rf_static_aad_length[968]       =   64'h0000000000000100;
assign   tb_i_aad[968]                        =   tb_i_aad[967];
assign   tb_i_rf_static_plaintext_length[968] =   64'h0000000000000280;
assign   tb_i_plaintext[968]                  =   tb_i_plaintext[967];
assign   tb_o_valid[968]                      =   1'b0;
assign   tb_o_sop[968]                        =   1'b0;
assign   tb_o_ciphertext[968]                 =   tb_o_ciphertext[967];
assign   tb_o_tag_ready[968]                  =   1'b0;
assign   tb_o_tag[968]                        =   tb_o_tag[967];

// CLK no. 969/1240
// *************************************************
assign   tb_i_valid[969]                      =   1'b0;
assign   tb_i_reset[969]                      =   1'b0;
assign   tb_i_sop[969]                        =   1'b0;
assign   tb_i_key_update[969]                 =   1'b0;
assign   tb_i_key[969]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[969]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[969]               =   1'b0;
assign   tb_i_rf_static_encrypt[969]          =   1'b1;
assign   tb_i_clear_fault_flags[969]          =   1'b0;
assign   tb_i_rf_static_aad_length[969]       =   64'h0000000000000100;
assign   tb_i_aad[969]                        =   tb_i_aad[968];
assign   tb_i_rf_static_plaintext_length[969] =   64'h0000000000000280;
assign   tb_i_plaintext[969]                  =   tb_i_plaintext[968];
assign   tb_o_valid[969]                      =   1'b0;
assign   tb_o_sop[969]                        =   1'b0;
assign   tb_o_ciphertext[969]                 =   tb_o_ciphertext[968];
assign   tb_o_tag_ready[969]                  =   1'b0;
assign   tb_o_tag[969]                        =   tb_o_tag[968];

// CLK no. 970/1240
// *************************************************
assign   tb_i_valid[970]                      =   1'b0;
assign   tb_i_reset[970]                      =   1'b0;
assign   tb_i_sop[970]                        =   1'b0;
assign   tb_i_key_update[970]                 =   1'b0;
assign   tb_i_key[970]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[970]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[970]               =   1'b0;
assign   tb_i_rf_static_encrypt[970]          =   1'b1;
assign   tb_i_clear_fault_flags[970]          =   1'b0;
assign   tb_i_rf_static_aad_length[970]       =   64'h0000000000000100;
assign   tb_i_aad[970]                        =   tb_i_aad[969];
assign   tb_i_rf_static_plaintext_length[970] =   64'h0000000000000280;
assign   tb_i_plaintext[970]                  =   tb_i_plaintext[969];
assign   tb_o_valid[970]                      =   1'b0;
assign   tb_o_sop[970]                        =   1'b0;
assign   tb_o_ciphertext[970]                 =   tb_o_ciphertext[969];
assign   tb_o_tag_ready[970]                  =   1'b0;
assign   tb_o_tag[970]                        =   tb_o_tag[969];

// CLK no. 971/1240
// *************************************************
assign   tb_i_valid[971]                      =   1'b0;
assign   tb_i_reset[971]                      =   1'b0;
assign   tb_i_sop[971]                        =   1'b0;
assign   tb_i_key_update[971]                 =   1'b0;
assign   tb_i_key[971]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[971]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[971]               =   1'b0;
assign   tb_i_rf_static_encrypt[971]          =   1'b1;
assign   tb_i_clear_fault_flags[971]          =   1'b0;
assign   tb_i_rf_static_aad_length[971]       =   64'h0000000000000100;
assign   tb_i_aad[971]                        =   tb_i_aad[970];
assign   tb_i_rf_static_plaintext_length[971] =   64'h0000000000000280;
assign   tb_i_plaintext[971]                  =   tb_i_plaintext[970];
assign   tb_o_valid[971]                      =   1'b0;
assign   tb_o_sop[971]                        =   1'b0;
assign   tb_o_ciphertext[971]                 =   tb_o_ciphertext[970];
assign   tb_o_tag_ready[971]                  =   1'b0;
assign   tb_o_tag[971]                        =   tb_o_tag[970];

// CLK no. 972/1240
// *************************************************
assign   tb_i_valid[972]                      =   1'b0;
assign   tb_i_reset[972]                      =   1'b0;
assign   tb_i_sop[972]                        =   1'b0;
assign   tb_i_key_update[972]                 =   1'b0;
assign   tb_i_key[972]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[972]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[972]               =   1'b0;
assign   tb_i_rf_static_encrypt[972]          =   1'b1;
assign   tb_i_clear_fault_flags[972]          =   1'b0;
assign   tb_i_rf_static_aad_length[972]       =   64'h0000000000000100;
assign   tb_i_aad[972]                        =   tb_i_aad[971];
assign   tb_i_rf_static_plaintext_length[972] =   64'h0000000000000280;
assign   tb_i_plaintext[972]                  =   tb_i_plaintext[971];
assign   tb_o_valid[972]                      =   1'b0;
assign   tb_o_sop[972]                        =   1'b0;
assign   tb_o_ciphertext[972]                 =   tb_o_ciphertext[971];
assign   tb_o_tag_ready[972]                  =   1'b0;
assign   tb_o_tag[972]                        =   tb_o_tag[971];

// CLK no. 973/1240
// *************************************************
assign   tb_i_valid[973]                      =   1'b0;
assign   tb_i_reset[973]                      =   1'b0;
assign   tb_i_sop[973]                        =   1'b0;
assign   tb_i_key_update[973]                 =   1'b0;
assign   tb_i_key[973]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[973]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[973]               =   1'b0;
assign   tb_i_rf_static_encrypt[973]          =   1'b1;
assign   tb_i_clear_fault_flags[973]          =   1'b0;
assign   tb_i_rf_static_aad_length[973]       =   64'h0000000000000100;
assign   tb_i_aad[973]                        =   tb_i_aad[972];
assign   tb_i_rf_static_plaintext_length[973] =   64'h0000000000000280;
assign   tb_i_plaintext[973]                  =   tb_i_plaintext[972];
assign   tb_o_valid[973]                      =   1'b0;
assign   tb_o_sop[973]                        =   1'b0;
assign   tb_o_ciphertext[973]                 =   tb_o_ciphertext[972];
assign   tb_o_tag_ready[973]                  =   1'b0;
assign   tb_o_tag[973]                        =   tb_o_tag[972];

// CLK no. 974/1240
// *************************************************
assign   tb_i_valid[974]                      =   1'b0;
assign   tb_i_reset[974]                      =   1'b0;
assign   tb_i_sop[974]                        =   1'b0;
assign   tb_i_key_update[974]                 =   1'b0;
assign   tb_i_key[974]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[974]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[974]               =   1'b0;
assign   tb_i_rf_static_encrypt[974]          =   1'b1;
assign   tb_i_clear_fault_flags[974]          =   1'b0;
assign   tb_i_rf_static_aad_length[974]       =   64'h0000000000000100;
assign   tb_i_aad[974]                        =   tb_i_aad[973];
assign   tb_i_rf_static_plaintext_length[974] =   64'h0000000000000280;
assign   tb_i_plaintext[974]                  =   tb_i_plaintext[973];
assign   tb_o_valid[974]                      =   1'b0;
assign   tb_o_sop[974]                        =   1'b0;
assign   tb_o_ciphertext[974]                 =   tb_o_ciphertext[973];
assign   tb_o_tag_ready[974]                  =   1'b0;
assign   tb_o_tag[974]                        =   tb_o_tag[973];

// CLK no. 975/1240
// *************************************************
assign   tb_i_valid[975]                      =   1'b0;
assign   tb_i_reset[975]                      =   1'b0;
assign   tb_i_sop[975]                        =   1'b0;
assign   tb_i_key_update[975]                 =   1'b0;
assign   tb_i_key[975]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[975]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[975]               =   1'b0;
assign   tb_i_rf_static_encrypt[975]          =   1'b1;
assign   tb_i_clear_fault_flags[975]          =   1'b0;
assign   tb_i_rf_static_aad_length[975]       =   64'h0000000000000100;
assign   tb_i_aad[975]                        =   tb_i_aad[974];
assign   tb_i_rf_static_plaintext_length[975] =   64'h0000000000000280;
assign   tb_i_plaintext[975]                  =   tb_i_plaintext[974];
assign   tb_o_valid[975]                      =   1'b0;
assign   tb_o_sop[975]                        =   1'b0;
assign   tb_o_ciphertext[975]                 =   tb_o_ciphertext[974];
assign   tb_o_tag_ready[975]                  =   1'b0;
assign   tb_o_tag[975]                        =   tb_o_tag[974];

// CLK no. 976/1240
// *************************************************
assign   tb_i_valid[976]                      =   1'b0;
assign   tb_i_reset[976]                      =   1'b0;
assign   tb_i_sop[976]                        =   1'b0;
assign   tb_i_key_update[976]                 =   1'b0;
assign   tb_i_key[976]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[976]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[976]               =   1'b0;
assign   tb_i_rf_static_encrypt[976]          =   1'b1;
assign   tb_i_clear_fault_flags[976]          =   1'b0;
assign   tb_i_rf_static_aad_length[976]       =   64'h0000000000000100;
assign   tb_i_aad[976]                        =   tb_i_aad[975];
assign   tb_i_rf_static_plaintext_length[976] =   64'h0000000000000280;
assign   tb_i_plaintext[976]                  =   tb_i_plaintext[975];
assign   tb_o_valid[976]                      =   1'b0;
assign   tb_o_sop[976]                        =   1'b0;
assign   tb_o_ciphertext[976]                 =   tb_o_ciphertext[975];
assign   tb_o_tag_ready[976]                  =   1'b0;
assign   tb_o_tag[976]                        =   tb_o_tag[975];

// CLK no. 977/1240
// *************************************************
assign   tb_i_valid[977]                      =   1'b0;
assign   tb_i_reset[977]                      =   1'b0;
assign   tb_i_sop[977]                        =   1'b0;
assign   tb_i_key_update[977]                 =   1'b0;
assign   tb_i_key[977]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[977]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[977]               =   1'b0;
assign   tb_i_rf_static_encrypt[977]          =   1'b1;
assign   tb_i_clear_fault_flags[977]          =   1'b0;
assign   tb_i_rf_static_aad_length[977]       =   64'h0000000000000100;
assign   tb_i_aad[977]                        =   tb_i_aad[976];
assign   tb_i_rf_static_plaintext_length[977] =   64'h0000000000000280;
assign   tb_i_plaintext[977]                  =   tb_i_plaintext[976];
assign   tb_o_valid[977]                      =   1'b0;
assign   tb_o_sop[977]                        =   1'b0;
assign   tb_o_ciphertext[977]                 =   tb_o_ciphertext[976];
assign   tb_o_tag_ready[977]                  =   1'b0;
assign   tb_o_tag[977]                        =   tb_o_tag[976];

// CLK no. 978/1240
// *************************************************
assign   tb_i_valid[978]                      =   1'b0;
assign   tb_i_reset[978]                      =   1'b0;
assign   tb_i_sop[978]                        =   1'b0;
assign   tb_i_key_update[978]                 =   1'b0;
assign   tb_i_key[978]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[978]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[978]               =   1'b0;
assign   tb_i_rf_static_encrypt[978]          =   1'b1;
assign   tb_i_clear_fault_flags[978]          =   1'b0;
assign   tb_i_rf_static_aad_length[978]       =   64'h0000000000000100;
assign   tb_i_aad[978]                        =   tb_i_aad[977];
assign   tb_i_rf_static_plaintext_length[978] =   64'h0000000000000280;
assign   tb_i_plaintext[978]                  =   tb_i_plaintext[977];
assign   tb_o_valid[978]                      =   1'b0;
assign   tb_o_sop[978]                        =   1'b0;
assign   tb_o_ciphertext[978]                 =   tb_o_ciphertext[977];
assign   tb_o_tag_ready[978]                  =   1'b0;
assign   tb_o_tag[978]                        =   tb_o_tag[977];

// CLK no. 979/1240
// *************************************************
assign   tb_i_valid[979]                      =   1'b0;
assign   tb_i_reset[979]                      =   1'b0;
assign   tb_i_sop[979]                        =   1'b0;
assign   tb_i_key_update[979]                 =   1'b0;
assign   tb_i_key[979]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[979]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[979]               =   1'b0;
assign   tb_i_rf_static_encrypt[979]          =   1'b1;
assign   tb_i_clear_fault_flags[979]          =   1'b0;
assign   tb_i_rf_static_aad_length[979]       =   64'h0000000000000100;
assign   tb_i_aad[979]                        =   tb_i_aad[978];
assign   tb_i_rf_static_plaintext_length[979] =   64'h0000000000000280;
assign   tb_i_plaintext[979]                  =   tb_i_plaintext[978];
assign   tb_o_valid[979]                      =   1'b0;
assign   tb_o_sop[979]                        =   1'b0;
assign   tb_o_ciphertext[979]                 =   tb_o_ciphertext[978];
assign   tb_o_tag_ready[979]                  =   1'b0;
assign   tb_o_tag[979]                        =   tb_o_tag[978];

// CLK no. 980/1240
// *************************************************
assign   tb_i_valid[980]                      =   1'b0;
assign   tb_i_reset[980]                      =   1'b0;
assign   tb_i_sop[980]                        =   1'b0;
assign   tb_i_key_update[980]                 =   1'b0;
assign   tb_i_key[980]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[980]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[980]               =   1'b0;
assign   tb_i_rf_static_encrypt[980]          =   1'b1;
assign   tb_i_clear_fault_flags[980]          =   1'b0;
assign   tb_i_rf_static_aad_length[980]       =   64'h0000000000000100;
assign   tb_i_aad[980]                        =   tb_i_aad[979];
assign   tb_i_rf_static_plaintext_length[980] =   64'h0000000000000280;
assign   tb_i_plaintext[980]                  =   tb_i_plaintext[979];
assign   tb_o_valid[980]                      =   1'b0;
assign   tb_o_sop[980]                        =   1'b0;
assign   tb_o_ciphertext[980]                 =   tb_o_ciphertext[979];
assign   tb_o_tag_ready[980]                  =   1'b0;
assign   tb_o_tag[980]                        =   tb_o_tag[979];

// CLK no. 981/1240
// *************************************************
assign   tb_i_valid[981]                      =   1'b0;
assign   tb_i_reset[981]                      =   1'b0;
assign   tb_i_sop[981]                        =   1'b0;
assign   tb_i_key_update[981]                 =   1'b0;
assign   tb_i_key[981]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[981]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[981]               =   1'b0;
assign   tb_i_rf_static_encrypt[981]          =   1'b1;
assign   tb_i_clear_fault_flags[981]          =   1'b0;
assign   tb_i_rf_static_aad_length[981]       =   64'h0000000000000100;
assign   tb_i_aad[981]                        =   tb_i_aad[980];
assign   tb_i_rf_static_plaintext_length[981] =   64'h0000000000000280;
assign   tb_i_plaintext[981]                  =   tb_i_plaintext[980];
assign   tb_o_valid[981]                      =   1'b0;
assign   tb_o_sop[981]                        =   1'b0;
assign   tb_o_ciphertext[981]                 =   tb_o_ciphertext[980];
assign   tb_o_tag_ready[981]                  =   1'b0;
assign   tb_o_tag[981]                        =   tb_o_tag[980];

// CLK no. 982/1240
// *************************************************
assign   tb_i_valid[982]                      =   1'b0;
assign   tb_i_reset[982]                      =   1'b0;
assign   tb_i_sop[982]                        =   1'b0;
assign   tb_i_key_update[982]                 =   1'b0;
assign   tb_i_key[982]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[982]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[982]               =   1'b0;
assign   tb_i_rf_static_encrypt[982]          =   1'b1;
assign   tb_i_clear_fault_flags[982]          =   1'b0;
assign   tb_i_rf_static_aad_length[982]       =   64'h0000000000000100;
assign   tb_i_aad[982]                        =   tb_i_aad[981];
assign   tb_i_rf_static_plaintext_length[982] =   64'h0000000000000280;
assign   tb_i_plaintext[982]                  =   tb_i_plaintext[981];
assign   tb_o_valid[982]                      =   1'b0;
assign   tb_o_sop[982]                        =   1'b0;
assign   tb_o_ciphertext[982]                 =   tb_o_ciphertext[981];
assign   tb_o_tag_ready[982]                  =   1'b0;
assign   tb_o_tag[982]                        =   tb_o_tag[981];

// CLK no. 983/1240
// *************************************************
assign   tb_i_valid[983]                      =   1'b0;
assign   tb_i_reset[983]                      =   1'b0;
assign   tb_i_sop[983]                        =   1'b0;
assign   tb_i_key_update[983]                 =   1'b0;
assign   tb_i_key[983]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[983]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[983]               =   1'b0;
assign   tb_i_rf_static_encrypt[983]          =   1'b1;
assign   tb_i_clear_fault_flags[983]          =   1'b0;
assign   tb_i_rf_static_aad_length[983]       =   64'h0000000000000100;
assign   tb_i_aad[983]                        =   tb_i_aad[982];
assign   tb_i_rf_static_plaintext_length[983] =   64'h0000000000000280;
assign   tb_i_plaintext[983]                  =   tb_i_plaintext[982];
assign   tb_o_valid[983]                      =   1'b0;
assign   tb_o_sop[983]                        =   1'b0;
assign   tb_o_ciphertext[983]                 =   tb_o_ciphertext[982];
assign   tb_o_tag_ready[983]                  =   1'b0;
assign   tb_o_tag[983]                        =   tb_o_tag[982];

// CLK no. 984/1240
// *************************************************
assign   tb_i_valid[984]                      =   1'b0;
assign   tb_i_reset[984]                      =   1'b0;
assign   tb_i_sop[984]                        =   1'b0;
assign   tb_i_key_update[984]                 =   1'b0;
assign   tb_i_key[984]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[984]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[984]               =   1'b0;
assign   tb_i_rf_static_encrypt[984]          =   1'b1;
assign   tb_i_clear_fault_flags[984]          =   1'b0;
assign   tb_i_rf_static_aad_length[984]       =   64'h0000000000000100;
assign   tb_i_aad[984]                        =   tb_i_aad[983];
assign   tb_i_rf_static_plaintext_length[984] =   64'h0000000000000280;
assign   tb_i_plaintext[984]                  =   tb_i_plaintext[983];
assign   tb_o_valid[984]                      =   1'b0;
assign   tb_o_sop[984]                        =   1'b0;
assign   tb_o_ciphertext[984]                 =   tb_o_ciphertext[983];
assign   tb_o_tag_ready[984]                  =   1'b0;
assign   tb_o_tag[984]                        =   tb_o_tag[983];

// CLK no. 985/1240
// *************************************************
assign   tb_i_valid[985]                      =   1'b0;
assign   tb_i_reset[985]                      =   1'b0;
assign   tb_i_sop[985]                        =   1'b0;
assign   tb_i_key_update[985]                 =   1'b0;
assign   tb_i_key[985]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[985]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[985]               =   1'b0;
assign   tb_i_rf_static_encrypt[985]          =   1'b1;
assign   tb_i_clear_fault_flags[985]          =   1'b0;
assign   tb_i_rf_static_aad_length[985]       =   64'h0000000000000100;
assign   tb_i_aad[985]                        =   tb_i_aad[984];
assign   tb_i_rf_static_plaintext_length[985] =   64'h0000000000000280;
assign   tb_i_plaintext[985]                  =   tb_i_plaintext[984];
assign   tb_o_valid[985]                      =   1'b0;
assign   tb_o_sop[985]                        =   1'b0;
assign   tb_o_ciphertext[985]                 =   tb_o_ciphertext[984];
assign   tb_o_tag_ready[985]                  =   1'b0;
assign   tb_o_tag[985]                        =   tb_o_tag[984];

// CLK no. 986/1240
// *************************************************
assign   tb_i_valid[986]                      =   1'b0;
assign   tb_i_reset[986]                      =   1'b0;
assign   tb_i_sop[986]                        =   1'b0;
assign   tb_i_key_update[986]                 =   1'b0;
assign   tb_i_key[986]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[986]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[986]               =   1'b0;
assign   tb_i_rf_static_encrypt[986]          =   1'b1;
assign   tb_i_clear_fault_flags[986]          =   1'b0;
assign   tb_i_rf_static_aad_length[986]       =   64'h0000000000000100;
assign   tb_i_aad[986]                        =   tb_i_aad[985];
assign   tb_i_rf_static_plaintext_length[986] =   64'h0000000000000280;
assign   tb_i_plaintext[986]                  =   tb_i_plaintext[985];
assign   tb_o_valid[986]                      =   1'b0;
assign   tb_o_sop[986]                        =   1'b0;
assign   tb_o_ciphertext[986]                 =   tb_o_ciphertext[985];
assign   tb_o_tag_ready[986]                  =   1'b0;
assign   tb_o_tag[986]                        =   tb_o_tag[985];

// CLK no. 987/1240
// *************************************************
assign   tb_i_valid[987]                      =   1'b0;
assign   tb_i_reset[987]                      =   1'b0;
assign   tb_i_sop[987]                        =   1'b0;
assign   tb_i_key_update[987]                 =   1'b0;
assign   tb_i_key[987]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[987]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[987]               =   1'b0;
assign   tb_i_rf_static_encrypt[987]          =   1'b1;
assign   tb_i_clear_fault_flags[987]          =   1'b0;
assign   tb_i_rf_static_aad_length[987]       =   64'h0000000000000100;
assign   tb_i_aad[987]                        =   tb_i_aad[986];
assign   tb_i_rf_static_plaintext_length[987] =   64'h0000000000000280;
assign   tb_i_plaintext[987]                  =   tb_i_plaintext[986];
assign   tb_o_valid[987]                      =   1'b0;
assign   tb_o_sop[987]                        =   1'b0;
assign   tb_o_ciphertext[987]                 =   tb_o_ciphertext[986];
assign   tb_o_tag_ready[987]                  =   1'b0;
assign   tb_o_tag[987]                        =   tb_o_tag[986];

// CLK no. 988/1240
// *************************************************
assign   tb_i_valid[988]                      =   1'b0;
assign   tb_i_reset[988]                      =   1'b0;
assign   tb_i_sop[988]                        =   1'b0;
assign   tb_i_key_update[988]                 =   1'b0;
assign   tb_i_key[988]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[988]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[988]               =   1'b0;
assign   tb_i_rf_static_encrypt[988]          =   1'b1;
assign   tb_i_clear_fault_flags[988]          =   1'b0;
assign   tb_i_rf_static_aad_length[988]       =   64'h0000000000000100;
assign   tb_i_aad[988]                        =   tb_i_aad[987];
assign   tb_i_rf_static_plaintext_length[988] =   64'h0000000000000280;
assign   tb_i_plaintext[988]                  =   tb_i_plaintext[987];
assign   tb_o_valid[988]                      =   1'b0;
assign   tb_o_sop[988]                        =   1'b0;
assign   tb_o_ciphertext[988]                 =   tb_o_ciphertext[987];
assign   tb_o_tag_ready[988]                  =   1'b0;
assign   tb_o_tag[988]                        =   tb_o_tag[987];

// CLK no. 989/1240
// *************************************************
assign   tb_i_valid[989]                      =   1'b0;
assign   tb_i_reset[989]                      =   1'b0;
assign   tb_i_sop[989]                        =   1'b0;
assign   tb_i_key_update[989]                 =   1'b0;
assign   tb_i_key[989]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[989]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[989]               =   1'b0;
assign   tb_i_rf_static_encrypt[989]          =   1'b1;
assign   tb_i_clear_fault_flags[989]          =   1'b0;
assign   tb_i_rf_static_aad_length[989]       =   64'h0000000000000100;
assign   tb_i_aad[989]                        =   tb_i_aad[988];
assign   tb_i_rf_static_plaintext_length[989] =   64'h0000000000000280;
assign   tb_i_plaintext[989]                  =   tb_i_plaintext[988];
assign   tb_o_valid[989]                      =   1'b0;
assign   tb_o_sop[989]                        =   1'b0;
assign   tb_o_ciphertext[989]                 =   tb_o_ciphertext[988];
assign   tb_o_tag_ready[989]                  =   1'b0;
assign   tb_o_tag[989]                        =   tb_o_tag[988];

// CLK no. 990/1240
// *************************************************
assign   tb_i_valid[990]                      =   1'b0;
assign   tb_i_reset[990]                      =   1'b0;
assign   tb_i_sop[990]                        =   1'b0;
assign   tb_i_key_update[990]                 =   1'b0;
assign   tb_i_key[990]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[990]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[990]               =   1'b0;
assign   tb_i_rf_static_encrypt[990]          =   1'b1;
assign   tb_i_clear_fault_flags[990]          =   1'b0;
assign   tb_i_rf_static_aad_length[990]       =   64'h0000000000000100;
assign   tb_i_aad[990]                        =   tb_i_aad[989];
assign   tb_i_rf_static_plaintext_length[990] =   64'h0000000000000280;
assign   tb_i_plaintext[990]                  =   tb_i_plaintext[989];
assign   tb_o_valid[990]                      =   1'b0;
assign   tb_o_sop[990]                        =   1'b0;
assign   tb_o_ciphertext[990]                 =   tb_o_ciphertext[989];
assign   tb_o_tag_ready[990]                  =   1'b0;
assign   tb_o_tag[990]                        =   tb_o_tag[989];

// CLK no. 991/1240
// *************************************************
assign   tb_i_valid[991]                      =   1'b0;
assign   tb_i_reset[991]                      =   1'b0;
assign   tb_i_sop[991]                        =   1'b0;
assign   tb_i_key_update[991]                 =   1'b0;
assign   tb_i_key[991]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[991]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[991]               =   1'b0;
assign   tb_i_rf_static_encrypt[991]          =   1'b1;
assign   tb_i_clear_fault_flags[991]          =   1'b0;
assign   tb_i_rf_static_aad_length[991]       =   64'h0000000000000100;
assign   tb_i_aad[991]                        =   tb_i_aad[990];
assign   tb_i_rf_static_plaintext_length[991] =   64'h0000000000000280;
assign   tb_i_plaintext[991]                  =   tb_i_plaintext[990];
assign   tb_o_valid[991]                      =   1'b1;
assign   tb_o_sop[991]                        =   1'b1;
assign   tb_o_ciphertext[991]                 =   256'h489e7ce0b958c302ca1c9c987199a8c21bafdc219f77a863352d0efce152b048;
assign   tb_o_tag_ready[991]                  =   1'b0;
assign   tb_o_tag[991]                        =   tb_o_tag[990];

// CLK no. 992/1240
// *************************************************
assign   tb_i_valid[992]                      =   1'b0;
assign   tb_i_reset[992]                      =   1'b0;
assign   tb_i_sop[992]                        =   1'b0;
assign   tb_i_key_update[992]                 =   1'b0;
assign   tb_i_key[992]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[992]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[992]               =   1'b0;
assign   tb_i_rf_static_encrypt[992]          =   1'b1;
assign   tb_i_clear_fault_flags[992]          =   1'b0;
assign   tb_i_rf_static_aad_length[992]       =   64'h0000000000000100;
assign   tb_i_aad[992]                        =   tb_i_aad[991];
assign   tb_i_rf_static_plaintext_length[992] =   64'h0000000000000280;
assign   tb_i_plaintext[992]                  =   tb_i_plaintext[991];
assign   tb_o_valid[992]                      =   1'b1;
assign   tb_o_sop[992]                        =   1'b0;
assign   tb_o_ciphertext[992]                 =   256'h984a53528677f183ebfa05fadb600b81e1eee5b0590764cb69099ffc73e240bf;
assign   tb_o_tag_ready[992]                  =   1'b0;
assign   tb_o_tag[992]                        =   tb_o_tag[991];

// CLK no. 993/1240
// *************************************************
assign   tb_i_valid[993]                      =   1'b0;
assign   tb_i_reset[993]                      =   1'b0;
assign   tb_i_sop[993]                        =   1'b0;
assign   tb_i_key_update[993]                 =   1'b0;
assign   tb_i_key[993]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[993]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[993]               =   1'b0;
assign   tb_i_rf_static_encrypt[993]          =   1'b1;
assign   tb_i_clear_fault_flags[993]          =   1'b0;
assign   tb_i_rf_static_aad_length[993]       =   64'h0000000000000100;
assign   tb_i_aad[993]                        =   tb_i_aad[992];
assign   tb_i_rf_static_plaintext_length[993] =   64'h0000000000000280;
assign   tb_i_plaintext[993]                  =   tb_i_plaintext[992];
assign   tb_o_valid[993]                      =   1'b1;
assign   tb_o_sop[993]                        =   1'b0;
assign   tb_o_ciphertext[993]                 =   256'h2de40e52eefc223bfa1dc0d906fed8ab;
assign   tb_o_tag_ready[993]                  =   1'b0;
assign   tb_o_tag[993]                        =   tb_o_tag[992];

// CLK no. 994/1240
// *************************************************
assign   tb_i_valid[994]                      =   1'b0;
assign   tb_i_reset[994]                      =   1'b0;
assign   tb_i_sop[994]                        =   1'b0;
assign   tb_i_key_update[994]                 =   1'b0;
assign   tb_i_key[994]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[994]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[994]               =   1'b0;
assign   tb_i_rf_static_encrypt[994]          =   1'b1;
assign   tb_i_clear_fault_flags[994]          =   1'b0;
assign   tb_i_rf_static_aad_length[994]       =   64'h0000000000000100;
assign   tb_i_aad[994]                        =   tb_i_aad[993];
assign   tb_i_rf_static_plaintext_length[994] =   64'h0000000000000280;
assign   tb_i_plaintext[994]                  =   tb_i_plaintext[993];
assign   tb_o_valid[994]                      =   1'b0;
assign   tb_o_sop[994]                        =   1'b0;
assign   tb_o_ciphertext[994]                 =   tb_o_ciphertext[993];
assign   tb_o_tag_ready[994]                  =   1'b0;
assign   tb_o_tag[994]                        =   tb_o_tag[993];

// CLK no. 995/1240
// *************************************************
assign   tb_i_valid[995]                      =   1'b0;
assign   tb_i_reset[995]                      =   1'b0;
assign   tb_i_sop[995]                        =   1'b0;
assign   tb_i_key_update[995]                 =   1'b0;
assign   tb_i_key[995]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[995]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[995]               =   1'b0;
assign   tb_i_rf_static_encrypt[995]          =   1'b1;
assign   tb_i_clear_fault_flags[995]          =   1'b0;
assign   tb_i_rf_static_aad_length[995]       =   64'h0000000000000100;
assign   tb_i_aad[995]                        =   tb_i_aad[994];
assign   tb_i_rf_static_plaintext_length[995] =   64'h0000000000000280;
assign   tb_i_plaintext[995]                  =   tb_i_plaintext[994];
assign   tb_o_valid[995]                      =   1'b0;
assign   tb_o_sop[995]                        =   1'b0;
assign   tb_o_ciphertext[995]                 =   tb_o_ciphertext[994];
assign   tb_o_tag_ready[995]                  =   1'b0;
assign   tb_o_tag[995]                        =   tb_o_tag[994];

// CLK no. 996/1240
// *************************************************
assign   tb_i_valid[996]                      =   1'b0;
assign   tb_i_reset[996]                      =   1'b0;
assign   tb_i_sop[996]                        =   1'b0;
assign   tb_i_key_update[996]                 =   1'b0;
assign   tb_i_key[996]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[996]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[996]               =   1'b0;
assign   tb_i_rf_static_encrypt[996]          =   1'b1;
assign   tb_i_clear_fault_flags[996]          =   1'b0;
assign   tb_i_rf_static_aad_length[996]       =   64'h0000000000000100;
assign   tb_i_aad[996]                        =   tb_i_aad[995];
assign   tb_i_rf_static_plaintext_length[996] =   64'h0000000000000280;
assign   tb_i_plaintext[996]                  =   tb_i_plaintext[995];
assign   tb_o_valid[996]                      =   1'b0;
assign   tb_o_sop[996]                        =   1'b0;
assign   tb_o_ciphertext[996]                 =   tb_o_ciphertext[995];
assign   tb_o_tag_ready[996]                  =   1'b0;
assign   tb_o_tag[996]                        =   tb_o_tag[995];

// CLK no. 997/1240
// *************************************************
assign   tb_i_valid[997]                      =   1'b0;
assign   tb_i_reset[997]                      =   1'b0;
assign   tb_i_sop[997]                        =   1'b0;
assign   tb_i_key_update[997]                 =   1'b0;
assign   tb_i_key[997]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[997]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[997]               =   1'b0;
assign   tb_i_rf_static_encrypt[997]          =   1'b1;
assign   tb_i_clear_fault_flags[997]          =   1'b0;
assign   tb_i_rf_static_aad_length[997]       =   64'h0000000000000100;
assign   tb_i_aad[997]                        =   tb_i_aad[996];
assign   tb_i_rf_static_plaintext_length[997] =   64'h0000000000000280;
assign   tb_i_plaintext[997]                  =   tb_i_plaintext[996];
assign   tb_o_valid[997]                      =   1'b0;
assign   tb_o_sop[997]                        =   1'b0;
assign   tb_o_ciphertext[997]                 =   tb_o_ciphertext[996];
assign   tb_o_tag_ready[997]                  =   1'b0;
assign   tb_o_tag[997]                        =   tb_o_tag[996];

// CLK no. 998/1240
// *************************************************
assign   tb_i_valid[998]                      =   1'b0;
assign   tb_i_reset[998]                      =   1'b0;
assign   tb_i_sop[998]                        =   1'b0;
assign   tb_i_key_update[998]                 =   1'b0;
assign   tb_i_key[998]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[998]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[998]               =   1'b0;
assign   tb_i_rf_static_encrypt[998]          =   1'b1;
assign   tb_i_clear_fault_flags[998]          =   1'b0;
assign   tb_i_rf_static_aad_length[998]       =   64'h0000000000000100;
assign   tb_i_aad[998]                        =   tb_i_aad[997];
assign   tb_i_rf_static_plaintext_length[998] =   64'h0000000000000280;
assign   tb_i_plaintext[998]                  =   tb_i_plaintext[997];
assign   tb_o_valid[998]                      =   1'b0;
assign   tb_o_sop[998]                        =   1'b0;
assign   tb_o_ciphertext[998]                 =   tb_o_ciphertext[997];
assign   tb_o_tag_ready[998]                  =   1'b0;
assign   tb_o_tag[998]                        =   tb_o_tag[997];

// CLK no. 999/1240
// *************************************************
assign   tb_i_valid[999]                      =   1'b0;
assign   tb_i_reset[999]                      =   1'b0;
assign   tb_i_sop[999]                        =   1'b0;
assign   tb_i_key_update[999]                 =   1'b0;
assign   tb_i_key[999]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[999]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[999]               =   1'b0;
assign   tb_i_rf_static_encrypt[999]          =   1'b1;
assign   tb_i_clear_fault_flags[999]          =   1'b0;
assign   tb_i_rf_static_aad_length[999]       =   64'h0000000000000100;
assign   tb_i_aad[999]                        =   tb_i_aad[998];
assign   tb_i_rf_static_plaintext_length[999] =   64'h0000000000000280;
assign   tb_i_plaintext[999]                  =   tb_i_plaintext[998];
assign   tb_o_valid[999]                      =   1'b0;
assign   tb_o_sop[999]                        =   1'b0;
assign   tb_o_ciphertext[999]                 =   tb_o_ciphertext[998];
assign   tb_o_tag_ready[999]                  =   1'b0;
assign   tb_o_tag[999]                        =   tb_o_tag[998];

// CLK no. 1000/1240
// *************************************************
assign   tb_i_valid[1000]                      =   1'b0;
assign   tb_i_reset[1000]                      =   1'b0;
assign   tb_i_sop[1000]                        =   1'b0;
assign   tb_i_key_update[1000]                 =   1'b0;
assign   tb_i_key[1000]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1000]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1000]               =   1'b0;
assign   tb_i_rf_static_encrypt[1000]          =   1'b1;
assign   tb_i_clear_fault_flags[1000]          =   1'b0;
assign   tb_i_rf_static_aad_length[1000]       =   64'h0000000000000100;
assign   tb_i_aad[1000]                        =   tb_i_aad[999];
assign   tb_i_rf_static_plaintext_length[1000] =   64'h0000000000000280;
assign   tb_i_plaintext[1000]                  =   tb_i_plaintext[999];
assign   tb_o_valid[1000]                      =   1'b0;
assign   tb_o_sop[1000]                        =   1'b0;
assign   tb_o_ciphertext[1000]                 =   tb_o_ciphertext[999];
assign   tb_o_tag_ready[1000]                  =   1'b0;
assign   tb_o_tag[1000]                        =   tb_o_tag[999];

// CLK no. 1001/1240
// *************************************************
assign   tb_i_valid[1001]                      =   1'b0;
assign   tb_i_reset[1001]                      =   1'b0;
assign   tb_i_sop[1001]                        =   1'b0;
assign   tb_i_key_update[1001]                 =   1'b0;
assign   tb_i_key[1001]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1001]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1001]               =   1'b0;
assign   tb_i_rf_static_encrypt[1001]          =   1'b1;
assign   tb_i_clear_fault_flags[1001]          =   1'b0;
assign   tb_i_rf_static_aad_length[1001]       =   64'h0000000000000100;
assign   tb_i_aad[1001]                        =   tb_i_aad[1000];
assign   tb_i_rf_static_plaintext_length[1001] =   64'h0000000000000280;
assign   tb_i_plaintext[1001]                  =   tb_i_plaintext[1000];
assign   tb_o_valid[1001]                      =   1'b0;
assign   tb_o_sop[1001]                        =   1'b0;
assign   tb_o_ciphertext[1001]                 =   tb_o_ciphertext[1000];
assign   tb_o_tag_ready[1001]                  =   1'b1;
assign   tb_o_tag[1001]                        =   128'h68bff9f8dbd2f76123f4191da9b19c6c;

// CLK no. 1002/1240
// *************************************************
assign   tb_i_valid[1002]                      =   1'b0;
assign   tb_i_reset[1002]                      =   1'b0;
assign   tb_i_sop[1002]                        =   1'b0;
assign   tb_i_key_update[1002]                 =   1'b0;
assign   tb_i_key[1002]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1002]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1002]               =   1'b0;
assign   tb_i_rf_static_encrypt[1002]          =   1'b1;
assign   tb_i_clear_fault_flags[1002]          =   1'b0;
assign   tb_i_rf_static_aad_length[1002]       =   64'h0000000000000100;
assign   tb_i_aad[1002]                        =   tb_i_aad[1001];
assign   tb_i_rf_static_plaintext_length[1002] =   64'h0000000000000280;
assign   tb_i_plaintext[1002]                  =   tb_i_plaintext[1001];
assign   tb_o_valid[1002]                      =   1'b0;
assign   tb_o_sop[1002]                        =   1'b0;
assign   tb_o_ciphertext[1002]                 =   tb_o_ciphertext[1001];
assign   tb_o_tag_ready[1002]                  =   1'b0;
assign   tb_o_tag[1002]                        =   tb_o_tag[1001];

// CLK no. 1003/1240
// *************************************************
assign   tb_i_valid[1003]                      =   1'b0;
assign   tb_i_reset[1003]                      =   1'b0;
assign   tb_i_sop[1003]                        =   1'b0;
assign   tb_i_key_update[1003]                 =   1'b0;
assign   tb_i_key[1003]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1003]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1003]               =   1'b0;
assign   tb_i_rf_static_encrypt[1003]          =   1'b1;
assign   tb_i_clear_fault_flags[1003]          =   1'b0;
assign   tb_i_rf_static_aad_length[1003]       =   64'h0000000000000100;
assign   tb_i_aad[1003]                        =   tb_i_aad[1002];
assign   tb_i_rf_static_plaintext_length[1003] =   64'h0000000000000280;
assign   tb_i_plaintext[1003]                  =   tb_i_plaintext[1002];
assign   tb_o_valid[1003]                      =   1'b0;
assign   tb_o_sop[1003]                        =   1'b0;
assign   tb_o_ciphertext[1003]                 =   tb_o_ciphertext[1002];
assign   tb_o_tag_ready[1003]                  =   1'b0;
assign   tb_o_tag[1003]                        =   tb_o_tag[1002];

// CLK no. 1004/1240
// *************************************************
assign   tb_i_valid[1004]                      =   1'b0;
assign   tb_i_reset[1004]                      =   1'b0;
assign   tb_i_sop[1004]                        =   1'b1;
assign   tb_i_key_update[1004]                 =   1'b0;
assign   tb_i_key[1004]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1004]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1004]               =   1'b0;
assign   tb_i_rf_static_encrypt[1004]          =   1'b1;
assign   tb_i_clear_fault_flags[1004]          =   1'b0;
assign   tb_i_rf_static_aad_length[1004]       =   64'h0000000000000100;
assign   tb_i_aad[1004]                        =   tb_i_aad[1003];
assign   tb_i_rf_static_plaintext_length[1004] =   64'h0000000000000280;
assign   tb_i_plaintext[1004]                  =   tb_i_plaintext[1003];
assign   tb_o_valid[1004]                      =   1'b0;
assign   tb_o_sop[1004]                        =   1'b0;
assign   tb_o_ciphertext[1004]                 =   tb_o_ciphertext[1003];
assign   tb_o_tag_ready[1004]                  =   1'b0;
assign   tb_o_tag[1004]                        =   tb_o_tag[1003];

// CLK no. 1005/1240
// *************************************************
assign   tb_i_valid[1005]                      =   1'b1;
assign   tb_i_reset[1005]                      =   1'b0;
assign   tb_i_sop[1005]                        =   1'b0;
assign   tb_i_key_update[1005]                 =   1'b0;
assign   tb_i_key[1005]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1005]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1005]               =   1'b0;
assign   tb_i_rf_static_encrypt[1005]          =   1'b1;
assign   tb_i_clear_fault_flags[1005]          =   1'b0;
assign   tb_i_rf_static_aad_length[1005]       =   64'h0000000000000100;
assign   tb_i_aad[1005]                        =   256'h0ea1d3a7b9bafe2e59a8352dc8f77570dfd293392097561de7f05de022d2470a;
assign   tb_i_rf_static_plaintext_length[1005] =   64'h0000000000000280;
assign   tb_i_plaintext[1005]                  =   tb_i_plaintext[1004];
assign   tb_o_valid[1005]                      =   1'b0;
assign   tb_o_sop[1005]                        =   1'b0;
assign   tb_o_ciphertext[1005]                 =   tb_o_ciphertext[1004];
assign   tb_o_tag_ready[1005]                  =   1'b0;
assign   tb_o_tag[1005]                        =   tb_o_tag[1004];

// CLK no. 1006/1240
// *************************************************
assign   tb_i_valid[1006]                      =   1'b1;
assign   tb_i_reset[1006]                      =   1'b0;
assign   tb_i_sop[1006]                        =   1'b0;
assign   tb_i_key_update[1006]                 =   1'b0;
assign   tb_i_key[1006]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1006]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1006]               =   1'b0;
assign   tb_i_rf_static_encrypt[1006]          =   1'b1;
assign   tb_i_clear_fault_flags[1006]          =   1'b0;
assign   tb_i_rf_static_aad_length[1006]       =   64'h0000000000000100;
assign   tb_i_aad[1006]                        =   tb_i_aad[1005];
assign   tb_i_rf_static_plaintext_length[1006] =   64'h0000000000000280;
assign   tb_i_plaintext[1006]                  =   256'hebeb2ee4e5b6249d14e61f2620bc92139427a297c9d8fdbea869b27a1fe4120c;
assign   tb_o_valid[1006]                      =   1'b0;
assign   tb_o_sop[1006]                        =   1'b0;
assign   tb_o_ciphertext[1006]                 =   tb_o_ciphertext[1005];
assign   tb_o_tag_ready[1006]                  =   1'b0;
assign   tb_o_tag[1006]                        =   tb_o_tag[1005];

// CLK no. 1007/1240
// *************************************************
assign   tb_i_valid[1007]                      =   1'b1;
assign   tb_i_reset[1007]                      =   1'b0;
assign   tb_i_sop[1007]                        =   1'b0;
assign   tb_i_key_update[1007]                 =   1'b0;
assign   tb_i_key[1007]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1007]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1007]               =   1'b0;
assign   tb_i_rf_static_encrypt[1007]          =   1'b1;
assign   tb_i_clear_fault_flags[1007]          =   1'b0;
assign   tb_i_rf_static_aad_length[1007]       =   64'h0000000000000100;
assign   tb_i_aad[1007]                        =   tb_i_aad[1006];
assign   tb_i_rf_static_plaintext_length[1007] =   64'h0000000000000280;
assign   tb_i_plaintext[1007]                  =   256'hba99d3da0e781ee6ae5e7c073ccccce524b9f5268c86831c7e726b3d256f318d;
assign   tb_o_valid[1007]                      =   1'b0;
assign   tb_o_sop[1007]                        =   1'b0;
assign   tb_o_ciphertext[1007]                 =   tb_o_ciphertext[1006];
assign   tb_o_tag_ready[1007]                  =   1'b0;
assign   tb_o_tag[1007]                        =   tb_o_tag[1006];

// CLK no. 1008/1240
// *************************************************
assign   tb_i_valid[1008]                      =   1'b1;
assign   tb_i_reset[1008]                      =   1'b0;
assign   tb_i_sop[1008]                        =   1'b0;
assign   tb_i_key_update[1008]                 =   1'b0;
assign   tb_i_key[1008]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1008]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1008]               =   1'b0;
assign   tb_i_rf_static_encrypt[1008]          =   1'b1;
assign   tb_i_clear_fault_flags[1008]          =   1'b0;
assign   tb_i_rf_static_aad_length[1008]       =   64'h0000000000000100;
assign   tb_i_aad[1008]                        =   tb_i_aad[1007];
assign   tb_i_rf_static_plaintext_length[1008] =   64'h0000000000000280;
assign   tb_i_plaintext[1008]                  =   256'haba82572f71fa9de39fe2168cfa80c25;
assign   tb_o_valid[1008]                      =   1'b0;
assign   tb_o_sop[1008]                        =   1'b0;
assign   tb_o_ciphertext[1008]                 =   tb_o_ciphertext[1007];
assign   tb_o_tag_ready[1008]                  =   1'b0;
assign   tb_o_tag[1008]                        =   tb_o_tag[1007];

// CLK no. 1009/1240
// *************************************************
assign   tb_i_valid[1009]                      =   1'b0;
assign   tb_i_reset[1009]                      =   1'b0;
assign   tb_i_sop[1009]                        =   1'b0;
assign   tb_i_key_update[1009]                 =   1'b0;
assign   tb_i_key[1009]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1009]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1009]               =   1'b0;
assign   tb_i_rf_static_encrypt[1009]          =   1'b1;
assign   tb_i_clear_fault_flags[1009]          =   1'b0;
assign   tb_i_rf_static_aad_length[1009]       =   64'h0000000000000100;
assign   tb_i_aad[1009]                        =   tb_i_aad[1008];
assign   tb_i_rf_static_plaintext_length[1009] =   64'h0000000000000280;
assign   tb_i_plaintext[1009]                  =   tb_i_plaintext[1008];
assign   tb_o_valid[1009]                      =   1'b0;
assign   tb_o_sop[1009]                        =   1'b0;
assign   tb_o_ciphertext[1009]                 =   tb_o_ciphertext[1008];
assign   tb_o_tag_ready[1009]                  =   1'b0;
assign   tb_o_tag[1009]                        =   tb_o_tag[1008];

// CLK no. 1010/1240
// *************************************************
assign   tb_i_valid[1010]                      =   1'b0;
assign   tb_i_reset[1010]                      =   1'b0;
assign   tb_i_sop[1010]                        =   1'b0;
assign   tb_i_key_update[1010]                 =   1'b0;
assign   tb_i_key[1010]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1010]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1010]               =   1'b0;
assign   tb_i_rf_static_encrypt[1010]          =   1'b1;
assign   tb_i_clear_fault_flags[1010]          =   1'b0;
assign   tb_i_rf_static_aad_length[1010]       =   64'h0000000000000100;
assign   tb_i_aad[1010]                        =   tb_i_aad[1009];
assign   tb_i_rf_static_plaintext_length[1010] =   64'h0000000000000280;
assign   tb_i_plaintext[1010]                  =   tb_i_plaintext[1009];
assign   tb_o_valid[1010]                      =   1'b0;
assign   tb_o_sop[1010]                        =   1'b0;
assign   tb_o_ciphertext[1010]                 =   tb_o_ciphertext[1009];
assign   tb_o_tag_ready[1010]                  =   1'b0;
assign   tb_o_tag[1010]                        =   tb_o_tag[1009];

// CLK no. 1011/1240
// *************************************************
assign   tb_i_valid[1011]                      =   1'b0;
assign   tb_i_reset[1011]                      =   1'b0;
assign   tb_i_sop[1011]                        =   1'b0;
assign   tb_i_key_update[1011]                 =   1'b0;
assign   tb_i_key[1011]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1011]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1011]               =   1'b0;
assign   tb_i_rf_static_encrypt[1011]          =   1'b1;
assign   tb_i_clear_fault_flags[1011]          =   1'b0;
assign   tb_i_rf_static_aad_length[1011]       =   64'h0000000000000100;
assign   tb_i_aad[1011]                        =   tb_i_aad[1010];
assign   tb_i_rf_static_plaintext_length[1011] =   64'h0000000000000280;
assign   tb_i_plaintext[1011]                  =   tb_i_plaintext[1010];
assign   tb_o_valid[1011]                      =   1'b0;
assign   tb_o_sop[1011]                        =   1'b0;
assign   tb_o_ciphertext[1011]                 =   tb_o_ciphertext[1010];
assign   tb_o_tag_ready[1011]                  =   1'b0;
assign   tb_o_tag[1011]                        =   tb_o_tag[1010];

// CLK no. 1012/1240
// *************************************************
assign   tb_i_valid[1012]                      =   1'b0;
assign   tb_i_reset[1012]                      =   1'b0;
assign   tb_i_sop[1012]                        =   1'b0;
assign   tb_i_key_update[1012]                 =   1'b0;
assign   tb_i_key[1012]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1012]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1012]               =   1'b0;
assign   tb_i_rf_static_encrypt[1012]          =   1'b1;
assign   tb_i_clear_fault_flags[1012]          =   1'b0;
assign   tb_i_rf_static_aad_length[1012]       =   64'h0000000000000100;
assign   tb_i_aad[1012]                        =   tb_i_aad[1011];
assign   tb_i_rf_static_plaintext_length[1012] =   64'h0000000000000280;
assign   tb_i_plaintext[1012]                  =   tb_i_plaintext[1011];
assign   tb_o_valid[1012]                      =   1'b0;
assign   tb_o_sop[1012]                        =   1'b0;
assign   tb_o_ciphertext[1012]                 =   tb_o_ciphertext[1011];
assign   tb_o_tag_ready[1012]                  =   1'b0;
assign   tb_o_tag[1012]                        =   tb_o_tag[1011];

// CLK no. 1013/1240
// *************************************************
assign   tb_i_valid[1013]                      =   1'b0;
assign   tb_i_reset[1013]                      =   1'b0;
assign   tb_i_sop[1013]                        =   1'b0;
assign   tb_i_key_update[1013]                 =   1'b0;
assign   tb_i_key[1013]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1013]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1013]               =   1'b0;
assign   tb_i_rf_static_encrypt[1013]          =   1'b1;
assign   tb_i_clear_fault_flags[1013]          =   1'b0;
assign   tb_i_rf_static_aad_length[1013]       =   64'h0000000000000100;
assign   tb_i_aad[1013]                        =   tb_i_aad[1012];
assign   tb_i_rf_static_plaintext_length[1013] =   64'h0000000000000280;
assign   tb_i_plaintext[1013]                  =   tb_i_plaintext[1012];
assign   tb_o_valid[1013]                      =   1'b0;
assign   tb_o_sop[1013]                        =   1'b0;
assign   tb_o_ciphertext[1013]                 =   tb_o_ciphertext[1012];
assign   tb_o_tag_ready[1013]                  =   1'b0;
assign   tb_o_tag[1013]                        =   tb_o_tag[1012];

// CLK no. 1014/1240
// *************************************************
assign   tb_i_valid[1014]                      =   1'b0;
assign   tb_i_reset[1014]                      =   1'b0;
assign   tb_i_sop[1014]                        =   1'b0;
assign   tb_i_key_update[1014]                 =   1'b0;
assign   tb_i_key[1014]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1014]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1014]               =   1'b0;
assign   tb_i_rf_static_encrypt[1014]          =   1'b1;
assign   tb_i_clear_fault_flags[1014]          =   1'b0;
assign   tb_i_rf_static_aad_length[1014]       =   64'h0000000000000100;
assign   tb_i_aad[1014]                        =   tb_i_aad[1013];
assign   tb_i_rf_static_plaintext_length[1014] =   64'h0000000000000280;
assign   tb_i_plaintext[1014]                  =   tb_i_plaintext[1013];
assign   tb_o_valid[1014]                      =   1'b0;
assign   tb_o_sop[1014]                        =   1'b0;
assign   tb_o_ciphertext[1014]                 =   tb_o_ciphertext[1013];
assign   tb_o_tag_ready[1014]                  =   1'b0;
assign   tb_o_tag[1014]                        =   tb_o_tag[1013];

// CLK no. 1015/1240
// *************************************************
assign   tb_i_valid[1015]                      =   1'b0;
assign   tb_i_reset[1015]                      =   1'b0;
assign   tb_i_sop[1015]                        =   1'b0;
assign   tb_i_key_update[1015]                 =   1'b0;
assign   tb_i_key[1015]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1015]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1015]               =   1'b0;
assign   tb_i_rf_static_encrypt[1015]          =   1'b1;
assign   tb_i_clear_fault_flags[1015]          =   1'b0;
assign   tb_i_rf_static_aad_length[1015]       =   64'h0000000000000100;
assign   tb_i_aad[1015]                        =   tb_i_aad[1014];
assign   tb_i_rf_static_plaintext_length[1015] =   64'h0000000000000280;
assign   tb_i_plaintext[1015]                  =   tb_i_plaintext[1014];
assign   tb_o_valid[1015]                      =   1'b0;
assign   tb_o_sop[1015]                        =   1'b0;
assign   tb_o_ciphertext[1015]                 =   tb_o_ciphertext[1014];
assign   tb_o_tag_ready[1015]                  =   1'b0;
assign   tb_o_tag[1015]                        =   tb_o_tag[1014];

// CLK no. 1016/1240
// *************************************************
assign   tb_i_valid[1016]                      =   1'b0;
assign   tb_i_reset[1016]                      =   1'b0;
assign   tb_i_sop[1016]                        =   1'b0;
assign   tb_i_key_update[1016]                 =   1'b0;
assign   tb_i_key[1016]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1016]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1016]               =   1'b0;
assign   tb_i_rf_static_encrypt[1016]          =   1'b1;
assign   tb_i_clear_fault_flags[1016]          =   1'b0;
assign   tb_i_rf_static_aad_length[1016]       =   64'h0000000000000100;
assign   tb_i_aad[1016]                        =   tb_i_aad[1015];
assign   tb_i_rf_static_plaintext_length[1016] =   64'h0000000000000280;
assign   tb_i_plaintext[1016]                  =   tb_i_plaintext[1015];
assign   tb_o_valid[1016]                      =   1'b0;
assign   tb_o_sop[1016]                        =   1'b0;
assign   tb_o_ciphertext[1016]                 =   tb_o_ciphertext[1015];
assign   tb_o_tag_ready[1016]                  =   1'b0;
assign   tb_o_tag[1016]                        =   tb_o_tag[1015];

// CLK no. 1017/1240
// *************************************************
assign   tb_i_valid[1017]                      =   1'b0;
assign   tb_i_reset[1017]                      =   1'b0;
assign   tb_i_sop[1017]                        =   1'b0;
assign   tb_i_key_update[1017]                 =   1'b0;
assign   tb_i_key[1017]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1017]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1017]               =   1'b0;
assign   tb_i_rf_static_encrypt[1017]          =   1'b1;
assign   tb_i_clear_fault_flags[1017]          =   1'b0;
assign   tb_i_rf_static_aad_length[1017]       =   64'h0000000000000100;
assign   tb_i_aad[1017]                        =   tb_i_aad[1016];
assign   tb_i_rf_static_plaintext_length[1017] =   64'h0000000000000280;
assign   tb_i_plaintext[1017]                  =   tb_i_plaintext[1016];
assign   tb_o_valid[1017]                      =   1'b0;
assign   tb_o_sop[1017]                        =   1'b0;
assign   tb_o_ciphertext[1017]                 =   tb_o_ciphertext[1016];
assign   tb_o_tag_ready[1017]                  =   1'b0;
assign   tb_o_tag[1017]                        =   tb_o_tag[1016];

// CLK no. 1018/1240
// *************************************************
assign   tb_i_valid[1018]                      =   1'b0;
assign   tb_i_reset[1018]                      =   1'b0;
assign   tb_i_sop[1018]                        =   1'b0;
assign   tb_i_key_update[1018]                 =   1'b0;
assign   tb_i_key[1018]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1018]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1018]               =   1'b0;
assign   tb_i_rf_static_encrypt[1018]          =   1'b1;
assign   tb_i_clear_fault_flags[1018]          =   1'b0;
assign   tb_i_rf_static_aad_length[1018]       =   64'h0000000000000100;
assign   tb_i_aad[1018]                        =   tb_i_aad[1017];
assign   tb_i_rf_static_plaintext_length[1018] =   64'h0000000000000280;
assign   tb_i_plaintext[1018]                  =   tb_i_plaintext[1017];
assign   tb_o_valid[1018]                      =   1'b0;
assign   tb_o_sop[1018]                        =   1'b0;
assign   tb_o_ciphertext[1018]                 =   tb_o_ciphertext[1017];
assign   tb_o_tag_ready[1018]                  =   1'b0;
assign   tb_o_tag[1018]                        =   tb_o_tag[1017];

// CLK no. 1019/1240
// *************************************************
assign   tb_i_valid[1019]                      =   1'b0;
assign   tb_i_reset[1019]                      =   1'b0;
assign   tb_i_sop[1019]                        =   1'b0;
assign   tb_i_key_update[1019]                 =   1'b0;
assign   tb_i_key[1019]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1019]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1019]               =   1'b0;
assign   tb_i_rf_static_encrypt[1019]          =   1'b1;
assign   tb_i_clear_fault_flags[1019]          =   1'b0;
assign   tb_i_rf_static_aad_length[1019]       =   64'h0000000000000100;
assign   tb_i_aad[1019]                        =   tb_i_aad[1018];
assign   tb_i_rf_static_plaintext_length[1019] =   64'h0000000000000280;
assign   tb_i_plaintext[1019]                  =   tb_i_plaintext[1018];
assign   tb_o_valid[1019]                      =   1'b0;
assign   tb_o_sop[1019]                        =   1'b0;
assign   tb_o_ciphertext[1019]                 =   tb_o_ciphertext[1018];
assign   tb_o_tag_ready[1019]                  =   1'b0;
assign   tb_o_tag[1019]                        =   tb_o_tag[1018];

// CLK no. 1020/1240
// *************************************************
assign   tb_i_valid[1020]                      =   1'b0;
assign   tb_i_reset[1020]                      =   1'b0;
assign   tb_i_sop[1020]                        =   1'b0;
assign   tb_i_key_update[1020]                 =   1'b0;
assign   tb_i_key[1020]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1020]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1020]               =   1'b0;
assign   tb_i_rf_static_encrypt[1020]          =   1'b1;
assign   tb_i_clear_fault_flags[1020]          =   1'b0;
assign   tb_i_rf_static_aad_length[1020]       =   64'h0000000000000100;
assign   tb_i_aad[1020]                        =   tb_i_aad[1019];
assign   tb_i_rf_static_plaintext_length[1020] =   64'h0000000000000280;
assign   tb_i_plaintext[1020]                  =   tb_i_plaintext[1019];
assign   tb_o_valid[1020]                      =   1'b0;
assign   tb_o_sop[1020]                        =   1'b0;
assign   tb_o_ciphertext[1020]                 =   tb_o_ciphertext[1019];
assign   tb_o_tag_ready[1020]                  =   1'b0;
assign   tb_o_tag[1020]                        =   tb_o_tag[1019];

// CLK no. 1021/1240
// *************************************************
assign   tb_i_valid[1021]                      =   1'b0;
assign   tb_i_reset[1021]                      =   1'b0;
assign   tb_i_sop[1021]                        =   1'b0;
assign   tb_i_key_update[1021]                 =   1'b0;
assign   tb_i_key[1021]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1021]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1021]               =   1'b0;
assign   tb_i_rf_static_encrypt[1021]          =   1'b1;
assign   tb_i_clear_fault_flags[1021]          =   1'b0;
assign   tb_i_rf_static_aad_length[1021]       =   64'h0000000000000100;
assign   tb_i_aad[1021]                        =   tb_i_aad[1020];
assign   tb_i_rf_static_plaintext_length[1021] =   64'h0000000000000280;
assign   tb_i_plaintext[1021]                  =   tb_i_plaintext[1020];
assign   tb_o_valid[1021]                      =   1'b0;
assign   tb_o_sop[1021]                        =   1'b0;
assign   tb_o_ciphertext[1021]                 =   tb_o_ciphertext[1020];
assign   tb_o_tag_ready[1021]                  =   1'b0;
assign   tb_o_tag[1021]                        =   tb_o_tag[1020];

// CLK no. 1022/1240
// *************************************************
assign   tb_i_valid[1022]                      =   1'b0;
assign   tb_i_reset[1022]                      =   1'b0;
assign   tb_i_sop[1022]                        =   1'b0;
assign   tb_i_key_update[1022]                 =   1'b0;
assign   tb_i_key[1022]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1022]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1022]               =   1'b0;
assign   tb_i_rf_static_encrypt[1022]          =   1'b1;
assign   tb_i_clear_fault_flags[1022]          =   1'b0;
assign   tb_i_rf_static_aad_length[1022]       =   64'h0000000000000100;
assign   tb_i_aad[1022]                        =   tb_i_aad[1021];
assign   tb_i_rf_static_plaintext_length[1022] =   64'h0000000000000280;
assign   tb_i_plaintext[1022]                  =   tb_i_plaintext[1021];
assign   tb_o_valid[1022]                      =   1'b0;
assign   tb_o_sop[1022]                        =   1'b0;
assign   tb_o_ciphertext[1022]                 =   tb_o_ciphertext[1021];
assign   tb_o_tag_ready[1022]                  =   1'b0;
assign   tb_o_tag[1022]                        =   tb_o_tag[1021];

// CLK no. 1023/1240
// *************************************************
assign   tb_i_valid[1023]                      =   1'b0;
assign   tb_i_reset[1023]                      =   1'b0;
assign   tb_i_sop[1023]                        =   1'b0;
assign   tb_i_key_update[1023]                 =   1'b0;
assign   tb_i_key[1023]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1023]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1023]               =   1'b0;
assign   tb_i_rf_static_encrypt[1023]          =   1'b1;
assign   tb_i_clear_fault_flags[1023]          =   1'b0;
assign   tb_i_rf_static_aad_length[1023]       =   64'h0000000000000100;
assign   tb_i_aad[1023]                        =   tb_i_aad[1022];
assign   tb_i_rf_static_plaintext_length[1023] =   64'h0000000000000280;
assign   tb_i_plaintext[1023]                  =   tb_i_plaintext[1022];
assign   tb_o_valid[1023]                      =   1'b0;
assign   tb_o_sop[1023]                        =   1'b0;
assign   tb_o_ciphertext[1023]                 =   tb_o_ciphertext[1022];
assign   tb_o_tag_ready[1023]                  =   1'b0;
assign   tb_o_tag[1023]                        =   tb_o_tag[1022];

// CLK no. 1024/1240
// *************************************************
assign   tb_i_valid[1024]                      =   1'b0;
assign   tb_i_reset[1024]                      =   1'b0;
assign   tb_i_sop[1024]                        =   1'b0;
assign   tb_i_key_update[1024]                 =   1'b0;
assign   tb_i_key[1024]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1024]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1024]               =   1'b0;
assign   tb_i_rf_static_encrypt[1024]          =   1'b1;
assign   tb_i_clear_fault_flags[1024]          =   1'b0;
assign   tb_i_rf_static_aad_length[1024]       =   64'h0000000000000100;
assign   tb_i_aad[1024]                        =   tb_i_aad[1023];
assign   tb_i_rf_static_plaintext_length[1024] =   64'h0000000000000280;
assign   tb_i_plaintext[1024]                  =   tb_i_plaintext[1023];
assign   tb_o_valid[1024]                      =   1'b0;
assign   tb_o_sop[1024]                        =   1'b0;
assign   tb_o_ciphertext[1024]                 =   tb_o_ciphertext[1023];
assign   tb_o_tag_ready[1024]                  =   1'b0;
assign   tb_o_tag[1024]                        =   tb_o_tag[1023];

// CLK no. 1025/1240
// *************************************************
assign   tb_i_valid[1025]                      =   1'b0;
assign   tb_i_reset[1025]                      =   1'b0;
assign   tb_i_sop[1025]                        =   1'b0;
assign   tb_i_key_update[1025]                 =   1'b0;
assign   tb_i_key[1025]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1025]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1025]               =   1'b0;
assign   tb_i_rf_static_encrypt[1025]          =   1'b1;
assign   tb_i_clear_fault_flags[1025]          =   1'b0;
assign   tb_i_rf_static_aad_length[1025]       =   64'h0000000000000100;
assign   tb_i_aad[1025]                        =   tb_i_aad[1024];
assign   tb_i_rf_static_plaintext_length[1025] =   64'h0000000000000280;
assign   tb_i_plaintext[1025]                  =   tb_i_plaintext[1024];
assign   tb_o_valid[1025]                      =   1'b0;
assign   tb_o_sop[1025]                        =   1'b0;
assign   tb_o_ciphertext[1025]                 =   tb_o_ciphertext[1024];
assign   tb_o_tag_ready[1025]                  =   1'b0;
assign   tb_o_tag[1025]                        =   tb_o_tag[1024];

// CLK no. 1026/1240
// *************************************************
assign   tb_i_valid[1026]                      =   1'b0;
assign   tb_i_reset[1026]                      =   1'b0;
assign   tb_i_sop[1026]                        =   1'b0;
assign   tb_i_key_update[1026]                 =   1'b0;
assign   tb_i_key[1026]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1026]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1026]               =   1'b0;
assign   tb_i_rf_static_encrypt[1026]          =   1'b1;
assign   tb_i_clear_fault_flags[1026]          =   1'b0;
assign   tb_i_rf_static_aad_length[1026]       =   64'h0000000000000100;
assign   tb_i_aad[1026]                        =   tb_i_aad[1025];
assign   tb_i_rf_static_plaintext_length[1026] =   64'h0000000000000280;
assign   tb_i_plaintext[1026]                  =   tb_i_plaintext[1025];
assign   tb_o_valid[1026]                      =   1'b0;
assign   tb_o_sop[1026]                        =   1'b0;
assign   tb_o_ciphertext[1026]                 =   tb_o_ciphertext[1025];
assign   tb_o_tag_ready[1026]                  =   1'b0;
assign   tb_o_tag[1026]                        =   tb_o_tag[1025];

// CLK no. 1027/1240
// *************************************************
assign   tb_i_valid[1027]                      =   1'b0;
assign   tb_i_reset[1027]                      =   1'b0;
assign   tb_i_sop[1027]                        =   1'b0;
assign   tb_i_key_update[1027]                 =   1'b0;
assign   tb_i_key[1027]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1027]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1027]               =   1'b0;
assign   tb_i_rf_static_encrypt[1027]          =   1'b1;
assign   tb_i_clear_fault_flags[1027]          =   1'b0;
assign   tb_i_rf_static_aad_length[1027]       =   64'h0000000000000100;
assign   tb_i_aad[1027]                        =   tb_i_aad[1026];
assign   tb_i_rf_static_plaintext_length[1027] =   64'h0000000000000280;
assign   tb_i_plaintext[1027]                  =   tb_i_plaintext[1026];
assign   tb_o_valid[1027]                      =   1'b0;
assign   tb_o_sop[1027]                        =   1'b0;
assign   tb_o_ciphertext[1027]                 =   tb_o_ciphertext[1026];
assign   tb_o_tag_ready[1027]                  =   1'b0;
assign   tb_o_tag[1027]                        =   tb_o_tag[1026];

// CLK no. 1028/1240
// *************************************************
assign   tb_i_valid[1028]                      =   1'b0;
assign   tb_i_reset[1028]                      =   1'b0;
assign   tb_i_sop[1028]                        =   1'b0;
assign   tb_i_key_update[1028]                 =   1'b0;
assign   tb_i_key[1028]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1028]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1028]               =   1'b0;
assign   tb_i_rf_static_encrypt[1028]          =   1'b1;
assign   tb_i_clear_fault_flags[1028]          =   1'b0;
assign   tb_i_rf_static_aad_length[1028]       =   64'h0000000000000100;
assign   tb_i_aad[1028]                        =   tb_i_aad[1027];
assign   tb_i_rf_static_plaintext_length[1028] =   64'h0000000000000280;
assign   tb_i_plaintext[1028]                  =   tb_i_plaintext[1027];
assign   tb_o_valid[1028]                      =   1'b0;
assign   tb_o_sop[1028]                        =   1'b0;
assign   tb_o_ciphertext[1028]                 =   tb_o_ciphertext[1027];
assign   tb_o_tag_ready[1028]                  =   1'b0;
assign   tb_o_tag[1028]                        =   tb_o_tag[1027];

// CLK no. 1029/1240
// *************************************************
assign   tb_i_valid[1029]                      =   1'b0;
assign   tb_i_reset[1029]                      =   1'b0;
assign   tb_i_sop[1029]                        =   1'b0;
assign   tb_i_key_update[1029]                 =   1'b0;
assign   tb_i_key[1029]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1029]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1029]               =   1'b0;
assign   tb_i_rf_static_encrypt[1029]          =   1'b1;
assign   tb_i_clear_fault_flags[1029]          =   1'b0;
assign   tb_i_rf_static_aad_length[1029]       =   64'h0000000000000100;
assign   tb_i_aad[1029]                        =   tb_i_aad[1028];
assign   tb_i_rf_static_plaintext_length[1029] =   64'h0000000000000280;
assign   tb_i_plaintext[1029]                  =   tb_i_plaintext[1028];
assign   tb_o_valid[1029]                      =   1'b0;
assign   tb_o_sop[1029]                        =   1'b0;
assign   tb_o_ciphertext[1029]                 =   tb_o_ciphertext[1028];
assign   tb_o_tag_ready[1029]                  =   1'b0;
assign   tb_o_tag[1029]                        =   tb_o_tag[1028];

// CLK no. 1030/1240
// *************************************************
assign   tb_i_valid[1030]                      =   1'b0;
assign   tb_i_reset[1030]                      =   1'b0;
assign   tb_i_sop[1030]                        =   1'b0;
assign   tb_i_key_update[1030]                 =   1'b0;
assign   tb_i_key[1030]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1030]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1030]               =   1'b0;
assign   tb_i_rf_static_encrypt[1030]          =   1'b1;
assign   tb_i_clear_fault_flags[1030]          =   1'b0;
assign   tb_i_rf_static_aad_length[1030]       =   64'h0000000000000100;
assign   tb_i_aad[1030]                        =   tb_i_aad[1029];
assign   tb_i_rf_static_plaintext_length[1030] =   64'h0000000000000280;
assign   tb_i_plaintext[1030]                  =   tb_i_plaintext[1029];
assign   tb_o_valid[1030]                      =   1'b0;
assign   tb_o_sop[1030]                        =   1'b0;
assign   tb_o_ciphertext[1030]                 =   tb_o_ciphertext[1029];
assign   tb_o_tag_ready[1030]                  =   1'b0;
assign   tb_o_tag[1030]                        =   tb_o_tag[1029];

// CLK no. 1031/1240
// *************************************************
assign   tb_i_valid[1031]                      =   1'b0;
assign   tb_i_reset[1031]                      =   1'b0;
assign   tb_i_sop[1031]                        =   1'b0;
assign   tb_i_key_update[1031]                 =   1'b0;
assign   tb_i_key[1031]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1031]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1031]               =   1'b0;
assign   tb_i_rf_static_encrypt[1031]          =   1'b1;
assign   tb_i_clear_fault_flags[1031]          =   1'b0;
assign   tb_i_rf_static_aad_length[1031]       =   64'h0000000000000100;
assign   tb_i_aad[1031]                        =   tb_i_aad[1030];
assign   tb_i_rf_static_plaintext_length[1031] =   64'h0000000000000280;
assign   tb_i_plaintext[1031]                  =   tb_i_plaintext[1030];
assign   tb_o_valid[1031]                      =   1'b0;
assign   tb_o_sop[1031]                        =   1'b0;
assign   tb_o_ciphertext[1031]                 =   tb_o_ciphertext[1030];
assign   tb_o_tag_ready[1031]                  =   1'b0;
assign   tb_o_tag[1031]                        =   tb_o_tag[1030];

// CLK no. 1032/1240
// *************************************************
assign   tb_i_valid[1032]                      =   1'b0;
assign   tb_i_reset[1032]                      =   1'b0;
assign   tb_i_sop[1032]                        =   1'b0;
assign   tb_i_key_update[1032]                 =   1'b0;
assign   tb_i_key[1032]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1032]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1032]               =   1'b0;
assign   tb_i_rf_static_encrypt[1032]          =   1'b1;
assign   tb_i_clear_fault_flags[1032]          =   1'b0;
assign   tb_i_rf_static_aad_length[1032]       =   64'h0000000000000100;
assign   tb_i_aad[1032]                        =   tb_i_aad[1031];
assign   tb_i_rf_static_plaintext_length[1032] =   64'h0000000000000280;
assign   tb_i_plaintext[1032]                  =   tb_i_plaintext[1031];
assign   tb_o_valid[1032]                      =   1'b0;
assign   tb_o_sop[1032]                        =   1'b0;
assign   tb_o_ciphertext[1032]                 =   tb_o_ciphertext[1031];
assign   tb_o_tag_ready[1032]                  =   1'b0;
assign   tb_o_tag[1032]                        =   tb_o_tag[1031];

// CLK no. 1033/1240
// *************************************************
assign   tb_i_valid[1033]                      =   1'b0;
assign   tb_i_reset[1033]                      =   1'b0;
assign   tb_i_sop[1033]                        =   1'b0;
assign   tb_i_key_update[1033]                 =   1'b0;
assign   tb_i_key[1033]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1033]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1033]               =   1'b0;
assign   tb_i_rf_static_encrypt[1033]          =   1'b1;
assign   tb_i_clear_fault_flags[1033]          =   1'b0;
assign   tb_i_rf_static_aad_length[1033]       =   64'h0000000000000100;
assign   tb_i_aad[1033]                        =   tb_i_aad[1032];
assign   tb_i_rf_static_plaintext_length[1033] =   64'h0000000000000280;
assign   tb_i_plaintext[1033]                  =   tb_i_plaintext[1032];
assign   tb_o_valid[1033]                      =   1'b0;
assign   tb_o_sop[1033]                        =   1'b0;
assign   tb_o_ciphertext[1033]                 =   tb_o_ciphertext[1032];
assign   tb_o_tag_ready[1033]                  =   1'b0;
assign   tb_o_tag[1033]                        =   tb_o_tag[1032];

// CLK no. 1034/1240
// *************************************************
assign   tb_i_valid[1034]                      =   1'b0;
assign   tb_i_reset[1034]                      =   1'b0;
assign   tb_i_sop[1034]                        =   1'b0;
assign   tb_i_key_update[1034]                 =   1'b0;
assign   tb_i_key[1034]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1034]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1034]               =   1'b0;
assign   tb_i_rf_static_encrypt[1034]          =   1'b1;
assign   tb_i_clear_fault_flags[1034]          =   1'b0;
assign   tb_i_rf_static_aad_length[1034]       =   64'h0000000000000100;
assign   tb_i_aad[1034]                        =   tb_i_aad[1033];
assign   tb_i_rf_static_plaintext_length[1034] =   64'h0000000000000280;
assign   tb_i_plaintext[1034]                  =   tb_i_plaintext[1033];
assign   tb_o_valid[1034]                      =   1'b0;
assign   tb_o_sop[1034]                        =   1'b0;
assign   tb_o_ciphertext[1034]                 =   tb_o_ciphertext[1033];
assign   tb_o_tag_ready[1034]                  =   1'b0;
assign   tb_o_tag[1034]                        =   tb_o_tag[1033];

// CLK no. 1035/1240
// *************************************************
assign   tb_i_valid[1035]                      =   1'b0;
assign   tb_i_reset[1035]                      =   1'b0;
assign   tb_i_sop[1035]                        =   1'b0;
assign   tb_i_key_update[1035]                 =   1'b0;
assign   tb_i_key[1035]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1035]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1035]               =   1'b0;
assign   tb_i_rf_static_encrypt[1035]          =   1'b1;
assign   tb_i_clear_fault_flags[1035]          =   1'b0;
assign   tb_i_rf_static_aad_length[1035]       =   64'h0000000000000100;
assign   tb_i_aad[1035]                        =   tb_i_aad[1034];
assign   tb_i_rf_static_plaintext_length[1035] =   64'h0000000000000280;
assign   tb_i_plaintext[1035]                  =   tb_i_plaintext[1034];
assign   tb_o_valid[1035]                      =   1'b0;
assign   tb_o_sop[1035]                        =   1'b0;
assign   tb_o_ciphertext[1035]                 =   tb_o_ciphertext[1034];
assign   tb_o_tag_ready[1035]                  =   1'b0;
assign   tb_o_tag[1035]                        =   tb_o_tag[1034];

// CLK no. 1036/1240
// *************************************************
assign   tb_i_valid[1036]                      =   1'b0;
assign   tb_i_reset[1036]                      =   1'b0;
assign   tb_i_sop[1036]                        =   1'b0;
assign   tb_i_key_update[1036]                 =   1'b0;
assign   tb_i_key[1036]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1036]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1036]               =   1'b0;
assign   tb_i_rf_static_encrypt[1036]          =   1'b1;
assign   tb_i_clear_fault_flags[1036]          =   1'b0;
assign   tb_i_rf_static_aad_length[1036]       =   64'h0000000000000100;
assign   tb_i_aad[1036]                        =   tb_i_aad[1035];
assign   tb_i_rf_static_plaintext_length[1036] =   64'h0000000000000280;
assign   tb_i_plaintext[1036]                  =   tb_i_plaintext[1035];
assign   tb_o_valid[1036]                      =   1'b0;
assign   tb_o_sop[1036]                        =   1'b0;
assign   tb_o_ciphertext[1036]                 =   tb_o_ciphertext[1035];
assign   tb_o_tag_ready[1036]                  =   1'b0;
assign   tb_o_tag[1036]                        =   tb_o_tag[1035];

// CLK no. 1037/1240
// *************************************************
assign   tb_i_valid[1037]                      =   1'b0;
assign   tb_i_reset[1037]                      =   1'b0;
assign   tb_i_sop[1037]                        =   1'b0;
assign   tb_i_key_update[1037]                 =   1'b0;
assign   tb_i_key[1037]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1037]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1037]               =   1'b0;
assign   tb_i_rf_static_encrypt[1037]          =   1'b1;
assign   tb_i_clear_fault_flags[1037]          =   1'b0;
assign   tb_i_rf_static_aad_length[1037]       =   64'h0000000000000100;
assign   tb_i_aad[1037]                        =   tb_i_aad[1036];
assign   tb_i_rf_static_plaintext_length[1037] =   64'h0000000000000280;
assign   tb_i_plaintext[1037]                  =   tb_i_plaintext[1036];
assign   tb_o_valid[1037]                      =   1'b0;
assign   tb_o_sop[1037]                        =   1'b0;
assign   tb_o_ciphertext[1037]                 =   tb_o_ciphertext[1036];
assign   tb_o_tag_ready[1037]                  =   1'b0;
assign   tb_o_tag[1037]                        =   tb_o_tag[1036];

// CLK no. 1038/1240
// *************************************************
assign   tb_i_valid[1038]                      =   1'b0;
assign   tb_i_reset[1038]                      =   1'b0;
assign   tb_i_sop[1038]                        =   1'b0;
assign   tb_i_key_update[1038]                 =   1'b0;
assign   tb_i_key[1038]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1038]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1038]               =   1'b0;
assign   tb_i_rf_static_encrypt[1038]          =   1'b1;
assign   tb_i_clear_fault_flags[1038]          =   1'b0;
assign   tb_i_rf_static_aad_length[1038]       =   64'h0000000000000100;
assign   tb_i_aad[1038]                        =   tb_i_aad[1037];
assign   tb_i_rf_static_plaintext_length[1038] =   64'h0000000000000280;
assign   tb_i_plaintext[1038]                  =   tb_i_plaintext[1037];
assign   tb_o_valid[1038]                      =   1'b0;
assign   tb_o_sop[1038]                        =   1'b0;
assign   tb_o_ciphertext[1038]                 =   tb_o_ciphertext[1037];
assign   tb_o_tag_ready[1038]                  =   1'b0;
assign   tb_o_tag[1038]                        =   tb_o_tag[1037];

// CLK no. 1039/1240
// *************************************************
assign   tb_i_valid[1039]                      =   1'b0;
assign   tb_i_reset[1039]                      =   1'b0;
assign   tb_i_sop[1039]                        =   1'b0;
assign   tb_i_key_update[1039]                 =   1'b0;
assign   tb_i_key[1039]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1039]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1039]               =   1'b0;
assign   tb_i_rf_static_encrypt[1039]          =   1'b1;
assign   tb_i_clear_fault_flags[1039]          =   1'b0;
assign   tb_i_rf_static_aad_length[1039]       =   64'h0000000000000100;
assign   tb_i_aad[1039]                        =   tb_i_aad[1038];
assign   tb_i_rf_static_plaintext_length[1039] =   64'h0000000000000280;
assign   tb_i_plaintext[1039]                  =   tb_i_plaintext[1038];
assign   tb_o_valid[1039]                      =   1'b0;
assign   tb_o_sop[1039]                        =   1'b0;
assign   tb_o_ciphertext[1039]                 =   tb_o_ciphertext[1038];
assign   tb_o_tag_ready[1039]                  =   1'b0;
assign   tb_o_tag[1039]                        =   tb_o_tag[1038];

// CLK no. 1040/1240
// *************************************************
assign   tb_i_valid[1040]                      =   1'b0;
assign   tb_i_reset[1040]                      =   1'b0;
assign   tb_i_sop[1040]                        =   1'b0;
assign   tb_i_key_update[1040]                 =   1'b0;
assign   tb_i_key[1040]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1040]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1040]               =   1'b0;
assign   tb_i_rf_static_encrypt[1040]          =   1'b1;
assign   tb_i_clear_fault_flags[1040]          =   1'b0;
assign   tb_i_rf_static_aad_length[1040]       =   64'h0000000000000100;
assign   tb_i_aad[1040]                        =   tb_i_aad[1039];
assign   tb_i_rf_static_plaintext_length[1040] =   64'h0000000000000280;
assign   tb_i_plaintext[1040]                  =   tb_i_plaintext[1039];
assign   tb_o_valid[1040]                      =   1'b0;
assign   tb_o_sop[1040]                        =   1'b0;
assign   tb_o_ciphertext[1040]                 =   tb_o_ciphertext[1039];
assign   tb_o_tag_ready[1040]                  =   1'b0;
assign   tb_o_tag[1040]                        =   tb_o_tag[1039];

// CLK no. 1041/1240
// *************************************************
assign   tb_i_valid[1041]                      =   1'b0;
assign   tb_i_reset[1041]                      =   1'b0;
assign   tb_i_sop[1041]                        =   1'b0;
assign   tb_i_key_update[1041]                 =   1'b0;
assign   tb_i_key[1041]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1041]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1041]               =   1'b0;
assign   tb_i_rf_static_encrypt[1041]          =   1'b1;
assign   tb_i_clear_fault_flags[1041]          =   1'b0;
assign   tb_i_rf_static_aad_length[1041]       =   64'h0000000000000100;
assign   tb_i_aad[1041]                        =   tb_i_aad[1040];
assign   tb_i_rf_static_plaintext_length[1041] =   64'h0000000000000280;
assign   tb_i_plaintext[1041]                  =   tb_i_plaintext[1040];
assign   tb_o_valid[1041]                      =   1'b0;
assign   tb_o_sop[1041]                        =   1'b0;
assign   tb_o_ciphertext[1041]                 =   tb_o_ciphertext[1040];
assign   tb_o_tag_ready[1041]                  =   1'b0;
assign   tb_o_tag[1041]                        =   tb_o_tag[1040];

// CLK no. 1042/1240
// *************************************************
assign   tb_i_valid[1042]                      =   1'b0;
assign   tb_i_reset[1042]                      =   1'b0;
assign   tb_i_sop[1042]                        =   1'b0;
assign   tb_i_key_update[1042]                 =   1'b0;
assign   tb_i_key[1042]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1042]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1042]               =   1'b0;
assign   tb_i_rf_static_encrypt[1042]          =   1'b1;
assign   tb_i_clear_fault_flags[1042]          =   1'b0;
assign   tb_i_rf_static_aad_length[1042]       =   64'h0000000000000100;
assign   tb_i_aad[1042]                        =   tb_i_aad[1041];
assign   tb_i_rf_static_plaintext_length[1042] =   64'h0000000000000280;
assign   tb_i_plaintext[1042]                  =   tb_i_plaintext[1041];
assign   tb_o_valid[1042]                      =   1'b0;
assign   tb_o_sop[1042]                        =   1'b0;
assign   tb_o_ciphertext[1042]                 =   tb_o_ciphertext[1041];
assign   tb_o_tag_ready[1042]                  =   1'b0;
assign   tb_o_tag[1042]                        =   tb_o_tag[1041];

// CLK no. 1043/1240
// *************************************************
assign   tb_i_valid[1043]                      =   1'b0;
assign   tb_i_reset[1043]                      =   1'b0;
assign   tb_i_sop[1043]                        =   1'b0;
assign   tb_i_key_update[1043]                 =   1'b0;
assign   tb_i_key[1043]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1043]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1043]               =   1'b0;
assign   tb_i_rf_static_encrypt[1043]          =   1'b1;
assign   tb_i_clear_fault_flags[1043]          =   1'b0;
assign   tb_i_rf_static_aad_length[1043]       =   64'h0000000000000100;
assign   tb_i_aad[1043]                        =   tb_i_aad[1042];
assign   tb_i_rf_static_plaintext_length[1043] =   64'h0000000000000280;
assign   tb_i_plaintext[1043]                  =   tb_i_plaintext[1042];
assign   tb_o_valid[1043]                      =   1'b0;
assign   tb_o_sop[1043]                        =   1'b0;
assign   tb_o_ciphertext[1043]                 =   tb_o_ciphertext[1042];
assign   tb_o_tag_ready[1043]                  =   1'b0;
assign   tb_o_tag[1043]                        =   tb_o_tag[1042];

// CLK no. 1044/1240
// *************************************************
assign   tb_i_valid[1044]                      =   1'b0;
assign   tb_i_reset[1044]                      =   1'b0;
assign   tb_i_sop[1044]                        =   1'b0;
assign   tb_i_key_update[1044]                 =   1'b0;
assign   tb_i_key[1044]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1044]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1044]               =   1'b0;
assign   tb_i_rf_static_encrypt[1044]          =   1'b1;
assign   tb_i_clear_fault_flags[1044]          =   1'b0;
assign   tb_i_rf_static_aad_length[1044]       =   64'h0000000000000100;
assign   tb_i_aad[1044]                        =   tb_i_aad[1043];
assign   tb_i_rf_static_plaintext_length[1044] =   64'h0000000000000280;
assign   tb_i_plaintext[1044]                  =   tb_i_plaintext[1043];
assign   tb_o_valid[1044]                      =   1'b0;
assign   tb_o_sop[1044]                        =   1'b0;
assign   tb_o_ciphertext[1044]                 =   tb_o_ciphertext[1043];
assign   tb_o_tag_ready[1044]                  =   1'b0;
assign   tb_o_tag[1044]                        =   tb_o_tag[1043];

// CLK no. 1045/1240
// *************************************************
assign   tb_i_valid[1045]                      =   1'b0;
assign   tb_i_reset[1045]                      =   1'b0;
assign   tb_i_sop[1045]                        =   1'b0;
assign   tb_i_key_update[1045]                 =   1'b0;
assign   tb_i_key[1045]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1045]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1045]               =   1'b0;
assign   tb_i_rf_static_encrypt[1045]          =   1'b1;
assign   tb_i_clear_fault_flags[1045]          =   1'b0;
assign   tb_i_rf_static_aad_length[1045]       =   64'h0000000000000100;
assign   tb_i_aad[1045]                        =   tb_i_aad[1044];
assign   tb_i_rf_static_plaintext_length[1045] =   64'h0000000000000280;
assign   tb_i_plaintext[1045]                  =   tb_i_plaintext[1044];
assign   tb_o_valid[1045]                      =   1'b0;
assign   tb_o_sop[1045]                        =   1'b0;
assign   tb_o_ciphertext[1045]                 =   tb_o_ciphertext[1044];
assign   tb_o_tag_ready[1045]                  =   1'b0;
assign   tb_o_tag[1045]                        =   tb_o_tag[1044];

// CLK no. 1046/1240
// *************************************************
assign   tb_i_valid[1046]                      =   1'b0;
assign   tb_i_reset[1046]                      =   1'b0;
assign   tb_i_sop[1046]                        =   1'b0;
assign   tb_i_key_update[1046]                 =   1'b0;
assign   tb_i_key[1046]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1046]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1046]               =   1'b0;
assign   tb_i_rf_static_encrypt[1046]          =   1'b1;
assign   tb_i_clear_fault_flags[1046]          =   1'b0;
assign   tb_i_rf_static_aad_length[1046]       =   64'h0000000000000100;
assign   tb_i_aad[1046]                        =   tb_i_aad[1045];
assign   tb_i_rf_static_plaintext_length[1046] =   64'h0000000000000280;
assign   tb_i_plaintext[1046]                  =   tb_i_plaintext[1045];
assign   tb_o_valid[1046]                      =   1'b0;
assign   tb_o_sop[1046]                        =   1'b0;
assign   tb_o_ciphertext[1046]                 =   tb_o_ciphertext[1045];
assign   tb_o_tag_ready[1046]                  =   1'b0;
assign   tb_o_tag[1046]                        =   tb_o_tag[1045];

// CLK no. 1047/1240
// *************************************************
assign   tb_i_valid[1047]                      =   1'b0;
assign   tb_i_reset[1047]                      =   1'b0;
assign   tb_i_sop[1047]                        =   1'b0;
assign   tb_i_key_update[1047]                 =   1'b0;
assign   tb_i_key[1047]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1047]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1047]               =   1'b0;
assign   tb_i_rf_static_encrypt[1047]          =   1'b1;
assign   tb_i_clear_fault_flags[1047]          =   1'b0;
assign   tb_i_rf_static_aad_length[1047]       =   64'h0000000000000100;
assign   tb_i_aad[1047]                        =   tb_i_aad[1046];
assign   tb_i_rf_static_plaintext_length[1047] =   64'h0000000000000280;
assign   tb_i_plaintext[1047]                  =   tb_i_plaintext[1046];
assign   tb_o_valid[1047]                      =   1'b0;
assign   tb_o_sop[1047]                        =   1'b0;
assign   tb_o_ciphertext[1047]                 =   tb_o_ciphertext[1046];
assign   tb_o_tag_ready[1047]                  =   1'b0;
assign   tb_o_tag[1047]                        =   tb_o_tag[1046];

// CLK no. 1048/1240
// *************************************************
assign   tb_i_valid[1048]                      =   1'b0;
assign   tb_i_reset[1048]                      =   1'b0;
assign   tb_i_sop[1048]                        =   1'b0;
assign   tb_i_key_update[1048]                 =   1'b0;
assign   tb_i_key[1048]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1048]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1048]               =   1'b0;
assign   tb_i_rf_static_encrypt[1048]          =   1'b1;
assign   tb_i_clear_fault_flags[1048]          =   1'b0;
assign   tb_i_rf_static_aad_length[1048]       =   64'h0000000000000100;
assign   tb_i_aad[1048]                        =   tb_i_aad[1047];
assign   tb_i_rf_static_plaintext_length[1048] =   64'h0000000000000280;
assign   tb_i_plaintext[1048]                  =   tb_i_plaintext[1047];
assign   tb_o_valid[1048]                      =   1'b0;
assign   tb_o_sop[1048]                        =   1'b0;
assign   tb_o_ciphertext[1048]                 =   tb_o_ciphertext[1047];
assign   tb_o_tag_ready[1048]                  =   1'b0;
assign   tb_o_tag[1048]                        =   tb_o_tag[1047];

// CLK no. 1049/1240
// *************************************************
assign   tb_i_valid[1049]                      =   1'b0;
assign   tb_i_reset[1049]                      =   1'b0;
assign   tb_i_sop[1049]                        =   1'b0;
assign   tb_i_key_update[1049]                 =   1'b0;
assign   tb_i_key[1049]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1049]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1049]               =   1'b0;
assign   tb_i_rf_static_encrypt[1049]          =   1'b1;
assign   tb_i_clear_fault_flags[1049]          =   1'b0;
assign   tb_i_rf_static_aad_length[1049]       =   64'h0000000000000100;
assign   tb_i_aad[1049]                        =   tb_i_aad[1048];
assign   tb_i_rf_static_plaintext_length[1049] =   64'h0000000000000280;
assign   tb_i_plaintext[1049]                  =   tb_i_plaintext[1048];
assign   tb_o_valid[1049]                      =   1'b0;
assign   tb_o_sop[1049]                        =   1'b0;
assign   tb_o_ciphertext[1049]                 =   tb_o_ciphertext[1048];
assign   tb_o_tag_ready[1049]                  =   1'b0;
assign   tb_o_tag[1049]                        =   tb_o_tag[1048];

// CLK no. 1050/1240
// *************************************************
assign   tb_i_valid[1050]                      =   1'b0;
assign   tb_i_reset[1050]                      =   1'b0;
assign   tb_i_sop[1050]                        =   1'b0;
assign   tb_i_key_update[1050]                 =   1'b0;
assign   tb_i_key[1050]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1050]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1050]               =   1'b0;
assign   tb_i_rf_static_encrypt[1050]          =   1'b1;
assign   tb_i_clear_fault_flags[1050]          =   1'b0;
assign   tb_i_rf_static_aad_length[1050]       =   64'h0000000000000100;
assign   tb_i_aad[1050]                        =   tb_i_aad[1049];
assign   tb_i_rf_static_plaintext_length[1050] =   64'h0000000000000280;
assign   tb_i_plaintext[1050]                  =   tb_i_plaintext[1049];
assign   tb_o_valid[1050]                      =   1'b1;
assign   tb_o_sop[1050]                        =   1'b1;
assign   tb_o_ciphertext[1050]                 =   256'h09760b6b4f67138e4f328da68fd8c9cb1f3b5142a80a865cf94f8c1c9a9576eb;
assign   tb_o_tag_ready[1050]                  =   1'b0;
assign   tb_o_tag[1050]                        =   tb_o_tag[1049];

// CLK no. 1051/1240
// *************************************************
assign   tb_i_valid[1051]                      =   1'b0;
assign   tb_i_reset[1051]                      =   1'b0;
assign   tb_i_sop[1051]                        =   1'b0;
assign   tb_i_key_update[1051]                 =   1'b0;
assign   tb_i_key[1051]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1051]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1051]               =   1'b0;
assign   tb_i_rf_static_encrypt[1051]          =   1'b1;
assign   tb_i_clear_fault_flags[1051]          =   1'b0;
assign   tb_i_rf_static_aad_length[1051]       =   64'h0000000000000100;
assign   tb_i_aad[1051]                        =   tb_i_aad[1050];
assign   tb_i_rf_static_plaintext_length[1051] =   64'h0000000000000280;
assign   tb_i_plaintext[1051]                  =   tb_i_plaintext[1050];
assign   tb_o_valid[1051]                      =   1'b1;
assign   tb_o_sop[1051]                        =   1'b0;
assign   tb_o_ciphertext[1051]                 =   256'hce05204c37cf82bba8f4f15cafe30b1db43577fb40e33172f60dee093a4b0c90;
assign   tb_o_tag_ready[1051]                  =   1'b0;
assign   tb_o_tag[1051]                        =   tb_o_tag[1050];

// CLK no. 1052/1240
// *************************************************
assign   tb_i_valid[1052]                      =   1'b0;
assign   tb_i_reset[1052]                      =   1'b0;
assign   tb_i_sop[1052]                        =   1'b0;
assign   tb_i_key_update[1052]                 =   1'b0;
assign   tb_i_key[1052]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1052]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1052]               =   1'b0;
assign   tb_i_rf_static_encrypt[1052]          =   1'b1;
assign   tb_i_clear_fault_flags[1052]          =   1'b0;
assign   tb_i_rf_static_aad_length[1052]       =   64'h0000000000000100;
assign   tb_i_aad[1052]                        =   tb_i_aad[1051];
assign   tb_i_rf_static_plaintext_length[1052] =   64'h0000000000000280;
assign   tb_i_plaintext[1052]                  =   tb_i_plaintext[1051];
assign   tb_o_valid[1052]                      =   1'b1;
assign   tb_o_sop[1052]                        =   1'b0;
assign   tb_o_ciphertext[1052]                 =   256'hcf075e2417f2d494716baf753950ecca;
assign   tb_o_tag_ready[1052]                  =   1'b0;
assign   tb_o_tag[1052]                        =   tb_o_tag[1051];

// CLK no. 1053/1240
// *************************************************
assign   tb_i_valid[1053]                      =   1'b0;
assign   tb_i_reset[1053]                      =   1'b0;
assign   tb_i_sop[1053]                        =   1'b0;
assign   tb_i_key_update[1053]                 =   1'b0;
assign   tb_i_key[1053]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1053]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1053]               =   1'b0;
assign   tb_i_rf_static_encrypt[1053]          =   1'b1;
assign   tb_i_clear_fault_flags[1053]          =   1'b0;
assign   tb_i_rf_static_aad_length[1053]       =   64'h0000000000000100;
assign   tb_i_aad[1053]                        =   tb_i_aad[1052];
assign   tb_i_rf_static_plaintext_length[1053] =   64'h0000000000000280;
assign   tb_i_plaintext[1053]                  =   tb_i_plaintext[1052];
assign   tb_o_valid[1053]                      =   1'b0;
assign   tb_o_sop[1053]                        =   1'b0;
assign   tb_o_ciphertext[1053]                 =   tb_o_ciphertext[1052];
assign   tb_o_tag_ready[1053]                  =   1'b0;
assign   tb_o_tag[1053]                        =   tb_o_tag[1052];

// CLK no. 1054/1240
// *************************************************
assign   tb_i_valid[1054]                      =   1'b0;
assign   tb_i_reset[1054]                      =   1'b0;
assign   tb_i_sop[1054]                        =   1'b0;
assign   tb_i_key_update[1054]                 =   1'b0;
assign   tb_i_key[1054]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1054]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1054]               =   1'b0;
assign   tb_i_rf_static_encrypt[1054]          =   1'b1;
assign   tb_i_clear_fault_flags[1054]          =   1'b0;
assign   tb_i_rf_static_aad_length[1054]       =   64'h0000000000000100;
assign   tb_i_aad[1054]                        =   tb_i_aad[1053];
assign   tb_i_rf_static_plaintext_length[1054] =   64'h0000000000000280;
assign   tb_i_plaintext[1054]                  =   tb_i_plaintext[1053];
assign   tb_o_valid[1054]                      =   1'b0;
assign   tb_o_sop[1054]                        =   1'b0;
assign   tb_o_ciphertext[1054]                 =   tb_o_ciphertext[1053];
assign   tb_o_tag_ready[1054]                  =   1'b0;
assign   tb_o_tag[1054]                        =   tb_o_tag[1053];

// CLK no. 1055/1240
// *************************************************
assign   tb_i_valid[1055]                      =   1'b0;
assign   tb_i_reset[1055]                      =   1'b0;
assign   tb_i_sop[1055]                        =   1'b0;
assign   tb_i_key_update[1055]                 =   1'b0;
assign   tb_i_key[1055]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1055]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1055]               =   1'b0;
assign   tb_i_rf_static_encrypt[1055]          =   1'b1;
assign   tb_i_clear_fault_flags[1055]          =   1'b0;
assign   tb_i_rf_static_aad_length[1055]       =   64'h0000000000000100;
assign   tb_i_aad[1055]                        =   tb_i_aad[1054];
assign   tb_i_rf_static_plaintext_length[1055] =   64'h0000000000000280;
assign   tb_i_plaintext[1055]                  =   tb_i_plaintext[1054];
assign   tb_o_valid[1055]                      =   1'b0;
assign   tb_o_sop[1055]                        =   1'b0;
assign   tb_o_ciphertext[1055]                 =   tb_o_ciphertext[1054];
assign   tb_o_tag_ready[1055]                  =   1'b0;
assign   tb_o_tag[1055]                        =   tb_o_tag[1054];

// CLK no. 1056/1240
// *************************************************
assign   tb_i_valid[1056]                      =   1'b0;
assign   tb_i_reset[1056]                      =   1'b0;
assign   tb_i_sop[1056]                        =   1'b0;
assign   tb_i_key_update[1056]                 =   1'b0;
assign   tb_i_key[1056]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1056]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1056]               =   1'b0;
assign   tb_i_rf_static_encrypt[1056]          =   1'b1;
assign   tb_i_clear_fault_flags[1056]          =   1'b0;
assign   tb_i_rf_static_aad_length[1056]       =   64'h0000000000000100;
assign   tb_i_aad[1056]                        =   tb_i_aad[1055];
assign   tb_i_rf_static_plaintext_length[1056] =   64'h0000000000000280;
assign   tb_i_plaintext[1056]                  =   tb_i_plaintext[1055];
assign   tb_o_valid[1056]                      =   1'b0;
assign   tb_o_sop[1056]                        =   1'b0;
assign   tb_o_ciphertext[1056]                 =   tb_o_ciphertext[1055];
assign   tb_o_tag_ready[1056]                  =   1'b0;
assign   tb_o_tag[1056]                        =   tb_o_tag[1055];

// CLK no. 1057/1240
// *************************************************
assign   tb_i_valid[1057]                      =   1'b0;
assign   tb_i_reset[1057]                      =   1'b0;
assign   tb_i_sop[1057]                        =   1'b0;
assign   tb_i_key_update[1057]                 =   1'b0;
assign   tb_i_key[1057]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1057]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1057]               =   1'b0;
assign   tb_i_rf_static_encrypt[1057]          =   1'b1;
assign   tb_i_clear_fault_flags[1057]          =   1'b0;
assign   tb_i_rf_static_aad_length[1057]       =   64'h0000000000000100;
assign   tb_i_aad[1057]                        =   tb_i_aad[1056];
assign   tb_i_rf_static_plaintext_length[1057] =   64'h0000000000000280;
assign   tb_i_plaintext[1057]                  =   tb_i_plaintext[1056];
assign   tb_o_valid[1057]                      =   1'b0;
assign   tb_o_sop[1057]                        =   1'b0;
assign   tb_o_ciphertext[1057]                 =   tb_o_ciphertext[1056];
assign   tb_o_tag_ready[1057]                  =   1'b0;
assign   tb_o_tag[1057]                        =   tb_o_tag[1056];

// CLK no. 1058/1240
// *************************************************
assign   tb_i_valid[1058]                      =   1'b0;
assign   tb_i_reset[1058]                      =   1'b0;
assign   tb_i_sop[1058]                        =   1'b0;
assign   tb_i_key_update[1058]                 =   1'b0;
assign   tb_i_key[1058]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1058]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1058]               =   1'b0;
assign   tb_i_rf_static_encrypt[1058]          =   1'b1;
assign   tb_i_clear_fault_flags[1058]          =   1'b0;
assign   tb_i_rf_static_aad_length[1058]       =   64'h0000000000000100;
assign   tb_i_aad[1058]                        =   tb_i_aad[1057];
assign   tb_i_rf_static_plaintext_length[1058] =   64'h0000000000000280;
assign   tb_i_plaintext[1058]                  =   tb_i_plaintext[1057];
assign   tb_o_valid[1058]                      =   1'b0;
assign   tb_o_sop[1058]                        =   1'b0;
assign   tb_o_ciphertext[1058]                 =   tb_o_ciphertext[1057];
assign   tb_o_tag_ready[1058]                  =   1'b0;
assign   tb_o_tag[1058]                        =   tb_o_tag[1057];

// CLK no. 1059/1240
// *************************************************
assign   tb_i_valid[1059]                      =   1'b0;
assign   tb_i_reset[1059]                      =   1'b0;
assign   tb_i_sop[1059]                        =   1'b0;
assign   tb_i_key_update[1059]                 =   1'b0;
assign   tb_i_key[1059]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1059]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1059]               =   1'b0;
assign   tb_i_rf_static_encrypt[1059]          =   1'b1;
assign   tb_i_clear_fault_flags[1059]          =   1'b0;
assign   tb_i_rf_static_aad_length[1059]       =   64'h0000000000000100;
assign   tb_i_aad[1059]                        =   tb_i_aad[1058];
assign   tb_i_rf_static_plaintext_length[1059] =   64'h0000000000000280;
assign   tb_i_plaintext[1059]                  =   tb_i_plaintext[1058];
assign   tb_o_valid[1059]                      =   1'b0;
assign   tb_o_sop[1059]                        =   1'b0;
assign   tb_o_ciphertext[1059]                 =   tb_o_ciphertext[1058];
assign   tb_o_tag_ready[1059]                  =   1'b0;
assign   tb_o_tag[1059]                        =   tb_o_tag[1058];

// CLK no. 1060/1240
// *************************************************
assign   tb_i_valid[1060]                      =   1'b0;
assign   tb_i_reset[1060]                      =   1'b0;
assign   tb_i_sop[1060]                        =   1'b0;
assign   tb_i_key_update[1060]                 =   1'b0;
assign   tb_i_key[1060]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1060]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1060]               =   1'b0;
assign   tb_i_rf_static_encrypt[1060]          =   1'b1;
assign   tb_i_clear_fault_flags[1060]          =   1'b0;
assign   tb_i_rf_static_aad_length[1060]       =   64'h0000000000000100;
assign   tb_i_aad[1060]                        =   tb_i_aad[1059];
assign   tb_i_rf_static_plaintext_length[1060] =   64'h0000000000000280;
assign   tb_i_plaintext[1060]                  =   tb_i_plaintext[1059];
assign   tb_o_valid[1060]                      =   1'b0;
assign   tb_o_sop[1060]                        =   1'b0;
assign   tb_o_ciphertext[1060]                 =   tb_o_ciphertext[1059];
assign   tb_o_tag_ready[1060]                  =   1'b1;
assign   tb_o_tag[1060]                        =   128'h2d41ff36f18dd474d36d423a0c61ff4e;

// CLK no. 1061/1240
// *************************************************
assign   tb_i_valid[1061]                      =   1'b0;
assign   tb_i_reset[1061]                      =   1'b0;
assign   tb_i_sop[1061]                        =   1'b0;
assign   tb_i_key_update[1061]                 =   1'b0;
assign   tb_i_key[1061]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1061]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1061]               =   1'b0;
assign   tb_i_rf_static_encrypt[1061]          =   1'b1;
assign   tb_i_clear_fault_flags[1061]          =   1'b0;
assign   tb_i_rf_static_aad_length[1061]       =   64'h0000000000000100;
assign   tb_i_aad[1061]                        =   tb_i_aad[1060];
assign   tb_i_rf_static_plaintext_length[1061] =   64'h0000000000000280;
assign   tb_i_plaintext[1061]                  =   tb_i_plaintext[1060];
assign   tb_o_valid[1061]                      =   1'b0;
assign   tb_o_sop[1061]                        =   1'b0;
assign   tb_o_ciphertext[1061]                 =   tb_o_ciphertext[1060];
assign   tb_o_tag_ready[1061]                  =   1'b0;
assign   tb_o_tag[1061]                        =   tb_o_tag[1060];

// CLK no. 1062/1240
// *************************************************
assign   tb_i_valid[1062]                      =   1'b0;
assign   tb_i_reset[1062]                      =   1'b0;
assign   tb_i_sop[1062]                        =   1'b0;
assign   tb_i_key_update[1062]                 =   1'b0;
assign   tb_i_key[1062]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1062]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1062]               =   1'b0;
assign   tb_i_rf_static_encrypt[1062]          =   1'b1;
assign   tb_i_clear_fault_flags[1062]          =   1'b0;
assign   tb_i_rf_static_aad_length[1062]       =   64'h0000000000000100;
assign   tb_i_aad[1062]                        =   tb_i_aad[1061];
assign   tb_i_rf_static_plaintext_length[1062] =   64'h0000000000000280;
assign   tb_i_plaintext[1062]                  =   tb_i_plaintext[1061];
assign   tb_o_valid[1062]                      =   1'b0;
assign   tb_o_sop[1062]                        =   1'b0;
assign   tb_o_ciphertext[1062]                 =   tb_o_ciphertext[1061];
assign   tb_o_tag_ready[1062]                  =   1'b0;
assign   tb_o_tag[1062]                        =   tb_o_tag[1061];

// CLK no. 1063/1240
// *************************************************
assign   tb_i_valid[1063]                      =   1'b0;
assign   tb_i_reset[1063]                      =   1'b0;
assign   tb_i_sop[1063]                        =   1'b1;
assign   tb_i_key_update[1063]                 =   1'b0;
assign   tb_i_key[1063]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1063]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1063]               =   1'b0;
assign   tb_i_rf_static_encrypt[1063]          =   1'b1;
assign   tb_i_clear_fault_flags[1063]          =   1'b0;
assign   tb_i_rf_static_aad_length[1063]       =   64'h0000000000000100;
assign   tb_i_aad[1063]                        =   tb_i_aad[1062];
assign   tb_i_rf_static_plaintext_length[1063] =   64'h0000000000000280;
assign   tb_i_plaintext[1063]                  =   tb_i_plaintext[1062];
assign   tb_o_valid[1063]                      =   1'b0;
assign   tb_o_sop[1063]                        =   1'b0;
assign   tb_o_ciphertext[1063]                 =   tb_o_ciphertext[1062];
assign   tb_o_tag_ready[1063]                  =   1'b0;
assign   tb_o_tag[1063]                        =   tb_o_tag[1062];

// CLK no. 1064/1240
// *************************************************
assign   tb_i_valid[1064]                      =   1'b1;
assign   tb_i_reset[1064]                      =   1'b0;
assign   tb_i_sop[1064]                        =   1'b0;
assign   tb_i_key_update[1064]                 =   1'b0;
assign   tb_i_key[1064]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1064]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1064]               =   1'b0;
assign   tb_i_rf_static_encrypt[1064]          =   1'b1;
assign   tb_i_clear_fault_flags[1064]          =   1'b0;
assign   tb_i_rf_static_aad_length[1064]       =   64'h0000000000000100;
assign   tb_i_aad[1064]                        =   256'h47ade441f76153376b1d6a9deee37886806f80411ef75d53f463698110d903a5;
assign   tb_i_rf_static_plaintext_length[1064] =   64'h0000000000000280;
assign   tb_i_plaintext[1064]                  =   tb_i_plaintext[1063];
assign   tb_o_valid[1064]                      =   1'b0;
assign   tb_o_sop[1064]                        =   1'b0;
assign   tb_o_ciphertext[1064]                 =   tb_o_ciphertext[1063];
assign   tb_o_tag_ready[1064]                  =   1'b0;
assign   tb_o_tag[1064]                        =   tb_o_tag[1063];

// CLK no. 1065/1240
// *************************************************
assign   tb_i_valid[1065]                      =   1'b1;
assign   tb_i_reset[1065]                      =   1'b0;
assign   tb_i_sop[1065]                        =   1'b0;
assign   tb_i_key_update[1065]                 =   1'b0;
assign   tb_i_key[1065]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1065]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1065]               =   1'b0;
assign   tb_i_rf_static_encrypt[1065]          =   1'b1;
assign   tb_i_clear_fault_flags[1065]          =   1'b0;
assign   tb_i_rf_static_aad_length[1065]       =   64'h0000000000000100;
assign   tb_i_aad[1065]                        =   tb_i_aad[1064];
assign   tb_i_rf_static_plaintext_length[1065] =   64'h0000000000000280;
assign   tb_i_plaintext[1065]                  =   256'hfb85431db40efd5fae5d8446e4458e4f352f1707d59b4758c73a2fae4061e4e4;
assign   tb_o_valid[1065]                      =   1'b0;
assign   tb_o_sop[1065]                        =   1'b0;
assign   tb_o_ciphertext[1065]                 =   tb_o_ciphertext[1064];
assign   tb_o_tag_ready[1065]                  =   1'b0;
assign   tb_o_tag[1065]                        =   tb_o_tag[1064];

// CLK no. 1066/1240
// *************************************************
assign   tb_i_valid[1066]                      =   1'b1;
assign   tb_i_reset[1066]                      =   1'b0;
assign   tb_i_sop[1066]                        =   1'b0;
assign   tb_i_key_update[1066]                 =   1'b0;
assign   tb_i_key[1066]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1066]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1066]               =   1'b0;
assign   tb_i_rf_static_encrypt[1066]          =   1'b1;
assign   tb_i_clear_fault_flags[1066]          =   1'b0;
assign   tb_i_rf_static_aad_length[1066]       =   64'h0000000000000100;
assign   tb_i_aad[1066]                        =   tb_i_aad[1065];
assign   tb_i_rf_static_plaintext_length[1066] =   64'h0000000000000280;
assign   tb_i_plaintext[1066]                  =   256'h72618c3fd748f3f8a9a0cd598a0a7fe7099c3df016a15436e9d64ac5b4e4fd60;
assign   tb_o_valid[1066]                      =   1'b0;
assign   tb_o_sop[1066]                        =   1'b0;
assign   tb_o_ciphertext[1066]                 =   tb_o_ciphertext[1065];
assign   tb_o_tag_ready[1066]                  =   1'b0;
assign   tb_o_tag[1066]                        =   tb_o_tag[1065];

// CLK no. 1067/1240
// *************************************************
assign   tb_i_valid[1067]                      =   1'b1;
assign   tb_i_reset[1067]                      =   1'b0;
assign   tb_i_sop[1067]                        =   1'b0;
assign   tb_i_key_update[1067]                 =   1'b0;
assign   tb_i_key[1067]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1067]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1067]               =   1'b0;
assign   tb_i_rf_static_encrypt[1067]          =   1'b1;
assign   tb_i_clear_fault_flags[1067]          =   1'b0;
assign   tb_i_rf_static_aad_length[1067]       =   64'h0000000000000100;
assign   tb_i_aad[1067]                        =   tb_i_aad[1066];
assign   tb_i_rf_static_plaintext_length[1067] =   64'h0000000000000280;
assign   tb_i_plaintext[1067]                  =   256'hf5ea1fcef266709482d103914e0effc2;
assign   tb_o_valid[1067]                      =   1'b0;
assign   tb_o_sop[1067]                        =   1'b0;
assign   tb_o_ciphertext[1067]                 =   tb_o_ciphertext[1066];
assign   tb_o_tag_ready[1067]                  =   1'b0;
assign   tb_o_tag[1067]                        =   tb_o_tag[1066];

// CLK no. 1068/1240
// *************************************************
assign   tb_i_valid[1068]                      =   1'b0;
assign   tb_i_reset[1068]                      =   1'b0;
assign   tb_i_sop[1068]                        =   1'b0;
assign   tb_i_key_update[1068]                 =   1'b0;
assign   tb_i_key[1068]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1068]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1068]               =   1'b0;
assign   tb_i_rf_static_encrypt[1068]          =   1'b1;
assign   tb_i_clear_fault_flags[1068]          =   1'b0;
assign   tb_i_rf_static_aad_length[1068]       =   64'h0000000000000100;
assign   tb_i_aad[1068]                        =   tb_i_aad[1067];
assign   tb_i_rf_static_plaintext_length[1068] =   64'h0000000000000280;
assign   tb_i_plaintext[1068]                  =   tb_i_plaintext[1067];
assign   tb_o_valid[1068]                      =   1'b0;
assign   tb_o_sop[1068]                        =   1'b0;
assign   tb_o_ciphertext[1068]                 =   tb_o_ciphertext[1067];
assign   tb_o_tag_ready[1068]                  =   1'b0;
assign   tb_o_tag[1068]                        =   tb_o_tag[1067];

// CLK no. 1069/1240
// *************************************************
assign   tb_i_valid[1069]                      =   1'b0;
assign   tb_i_reset[1069]                      =   1'b0;
assign   tb_i_sop[1069]                        =   1'b0;
assign   tb_i_key_update[1069]                 =   1'b0;
assign   tb_i_key[1069]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1069]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1069]               =   1'b0;
assign   tb_i_rf_static_encrypt[1069]          =   1'b1;
assign   tb_i_clear_fault_flags[1069]          =   1'b0;
assign   tb_i_rf_static_aad_length[1069]       =   64'h0000000000000100;
assign   tb_i_aad[1069]                        =   tb_i_aad[1068];
assign   tb_i_rf_static_plaintext_length[1069] =   64'h0000000000000280;
assign   tb_i_plaintext[1069]                  =   tb_i_plaintext[1068];
assign   tb_o_valid[1069]                      =   1'b0;
assign   tb_o_sop[1069]                        =   1'b0;
assign   tb_o_ciphertext[1069]                 =   tb_o_ciphertext[1068];
assign   tb_o_tag_ready[1069]                  =   1'b0;
assign   tb_o_tag[1069]                        =   tb_o_tag[1068];

// CLK no. 1070/1240
// *************************************************
assign   tb_i_valid[1070]                      =   1'b0;
assign   tb_i_reset[1070]                      =   1'b0;
assign   tb_i_sop[1070]                        =   1'b0;
assign   tb_i_key_update[1070]                 =   1'b0;
assign   tb_i_key[1070]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1070]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1070]               =   1'b0;
assign   tb_i_rf_static_encrypt[1070]          =   1'b1;
assign   tb_i_clear_fault_flags[1070]          =   1'b0;
assign   tb_i_rf_static_aad_length[1070]       =   64'h0000000000000100;
assign   tb_i_aad[1070]                        =   tb_i_aad[1069];
assign   tb_i_rf_static_plaintext_length[1070] =   64'h0000000000000280;
assign   tb_i_plaintext[1070]                  =   tb_i_plaintext[1069];
assign   tb_o_valid[1070]                      =   1'b0;
assign   tb_o_sop[1070]                        =   1'b0;
assign   tb_o_ciphertext[1070]                 =   tb_o_ciphertext[1069];
assign   tb_o_tag_ready[1070]                  =   1'b0;
assign   tb_o_tag[1070]                        =   tb_o_tag[1069];

// CLK no. 1071/1240
// *************************************************
assign   tb_i_valid[1071]                      =   1'b0;
assign   tb_i_reset[1071]                      =   1'b0;
assign   tb_i_sop[1071]                        =   1'b0;
assign   tb_i_key_update[1071]                 =   1'b0;
assign   tb_i_key[1071]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1071]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1071]               =   1'b0;
assign   tb_i_rf_static_encrypt[1071]          =   1'b1;
assign   tb_i_clear_fault_flags[1071]          =   1'b0;
assign   tb_i_rf_static_aad_length[1071]       =   64'h0000000000000100;
assign   tb_i_aad[1071]                        =   tb_i_aad[1070];
assign   tb_i_rf_static_plaintext_length[1071] =   64'h0000000000000280;
assign   tb_i_plaintext[1071]                  =   tb_i_plaintext[1070];
assign   tb_o_valid[1071]                      =   1'b0;
assign   tb_o_sop[1071]                        =   1'b0;
assign   tb_o_ciphertext[1071]                 =   tb_o_ciphertext[1070];
assign   tb_o_tag_ready[1071]                  =   1'b0;
assign   tb_o_tag[1071]                        =   tb_o_tag[1070];

// CLK no. 1072/1240
// *************************************************
assign   tb_i_valid[1072]                      =   1'b0;
assign   tb_i_reset[1072]                      =   1'b0;
assign   tb_i_sop[1072]                        =   1'b0;
assign   tb_i_key_update[1072]                 =   1'b0;
assign   tb_i_key[1072]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1072]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1072]               =   1'b0;
assign   tb_i_rf_static_encrypt[1072]          =   1'b1;
assign   tb_i_clear_fault_flags[1072]          =   1'b0;
assign   tb_i_rf_static_aad_length[1072]       =   64'h0000000000000100;
assign   tb_i_aad[1072]                        =   tb_i_aad[1071];
assign   tb_i_rf_static_plaintext_length[1072] =   64'h0000000000000280;
assign   tb_i_plaintext[1072]                  =   tb_i_plaintext[1071];
assign   tb_o_valid[1072]                      =   1'b0;
assign   tb_o_sop[1072]                        =   1'b0;
assign   tb_o_ciphertext[1072]                 =   tb_o_ciphertext[1071];
assign   tb_o_tag_ready[1072]                  =   1'b0;
assign   tb_o_tag[1072]                        =   tb_o_tag[1071];

// CLK no. 1073/1240
// *************************************************
assign   tb_i_valid[1073]                      =   1'b0;
assign   tb_i_reset[1073]                      =   1'b0;
assign   tb_i_sop[1073]                        =   1'b0;
assign   tb_i_key_update[1073]                 =   1'b0;
assign   tb_i_key[1073]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1073]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1073]               =   1'b0;
assign   tb_i_rf_static_encrypt[1073]          =   1'b1;
assign   tb_i_clear_fault_flags[1073]          =   1'b0;
assign   tb_i_rf_static_aad_length[1073]       =   64'h0000000000000100;
assign   tb_i_aad[1073]                        =   tb_i_aad[1072];
assign   tb_i_rf_static_plaintext_length[1073] =   64'h0000000000000280;
assign   tb_i_plaintext[1073]                  =   tb_i_plaintext[1072];
assign   tb_o_valid[1073]                      =   1'b0;
assign   tb_o_sop[1073]                        =   1'b0;
assign   tb_o_ciphertext[1073]                 =   tb_o_ciphertext[1072];
assign   tb_o_tag_ready[1073]                  =   1'b0;
assign   tb_o_tag[1073]                        =   tb_o_tag[1072];

// CLK no. 1074/1240
// *************************************************
assign   tb_i_valid[1074]                      =   1'b0;
assign   tb_i_reset[1074]                      =   1'b0;
assign   tb_i_sop[1074]                        =   1'b0;
assign   tb_i_key_update[1074]                 =   1'b0;
assign   tb_i_key[1074]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1074]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1074]               =   1'b0;
assign   tb_i_rf_static_encrypt[1074]          =   1'b1;
assign   tb_i_clear_fault_flags[1074]          =   1'b0;
assign   tb_i_rf_static_aad_length[1074]       =   64'h0000000000000100;
assign   tb_i_aad[1074]                        =   tb_i_aad[1073];
assign   tb_i_rf_static_plaintext_length[1074] =   64'h0000000000000280;
assign   tb_i_plaintext[1074]                  =   tb_i_plaintext[1073];
assign   tb_o_valid[1074]                      =   1'b0;
assign   tb_o_sop[1074]                        =   1'b0;
assign   tb_o_ciphertext[1074]                 =   tb_o_ciphertext[1073];
assign   tb_o_tag_ready[1074]                  =   1'b0;
assign   tb_o_tag[1074]                        =   tb_o_tag[1073];

// CLK no. 1075/1240
// *************************************************
assign   tb_i_valid[1075]                      =   1'b0;
assign   tb_i_reset[1075]                      =   1'b0;
assign   tb_i_sop[1075]                        =   1'b0;
assign   tb_i_key_update[1075]                 =   1'b0;
assign   tb_i_key[1075]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1075]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1075]               =   1'b0;
assign   tb_i_rf_static_encrypt[1075]          =   1'b1;
assign   tb_i_clear_fault_flags[1075]          =   1'b0;
assign   tb_i_rf_static_aad_length[1075]       =   64'h0000000000000100;
assign   tb_i_aad[1075]                        =   tb_i_aad[1074];
assign   tb_i_rf_static_plaintext_length[1075] =   64'h0000000000000280;
assign   tb_i_plaintext[1075]                  =   tb_i_plaintext[1074];
assign   tb_o_valid[1075]                      =   1'b0;
assign   tb_o_sop[1075]                        =   1'b0;
assign   tb_o_ciphertext[1075]                 =   tb_o_ciphertext[1074];
assign   tb_o_tag_ready[1075]                  =   1'b0;
assign   tb_o_tag[1075]                        =   tb_o_tag[1074];

// CLK no. 1076/1240
// *************************************************
assign   tb_i_valid[1076]                      =   1'b0;
assign   tb_i_reset[1076]                      =   1'b0;
assign   tb_i_sop[1076]                        =   1'b0;
assign   tb_i_key_update[1076]                 =   1'b0;
assign   tb_i_key[1076]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1076]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1076]               =   1'b0;
assign   tb_i_rf_static_encrypt[1076]          =   1'b1;
assign   tb_i_clear_fault_flags[1076]          =   1'b0;
assign   tb_i_rf_static_aad_length[1076]       =   64'h0000000000000100;
assign   tb_i_aad[1076]                        =   tb_i_aad[1075];
assign   tb_i_rf_static_plaintext_length[1076] =   64'h0000000000000280;
assign   tb_i_plaintext[1076]                  =   tb_i_plaintext[1075];
assign   tb_o_valid[1076]                      =   1'b0;
assign   tb_o_sop[1076]                        =   1'b0;
assign   tb_o_ciphertext[1076]                 =   tb_o_ciphertext[1075];
assign   tb_o_tag_ready[1076]                  =   1'b0;
assign   tb_o_tag[1076]                        =   tb_o_tag[1075];

// CLK no. 1077/1240
// *************************************************
assign   tb_i_valid[1077]                      =   1'b0;
assign   tb_i_reset[1077]                      =   1'b0;
assign   tb_i_sop[1077]                        =   1'b0;
assign   tb_i_key_update[1077]                 =   1'b0;
assign   tb_i_key[1077]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1077]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1077]               =   1'b0;
assign   tb_i_rf_static_encrypt[1077]          =   1'b1;
assign   tb_i_clear_fault_flags[1077]          =   1'b0;
assign   tb_i_rf_static_aad_length[1077]       =   64'h0000000000000100;
assign   tb_i_aad[1077]                        =   tb_i_aad[1076];
assign   tb_i_rf_static_plaintext_length[1077] =   64'h0000000000000280;
assign   tb_i_plaintext[1077]                  =   tb_i_plaintext[1076];
assign   tb_o_valid[1077]                      =   1'b0;
assign   tb_o_sop[1077]                        =   1'b0;
assign   tb_o_ciphertext[1077]                 =   tb_o_ciphertext[1076];
assign   tb_o_tag_ready[1077]                  =   1'b0;
assign   tb_o_tag[1077]                        =   tb_o_tag[1076];

// CLK no. 1078/1240
// *************************************************
assign   tb_i_valid[1078]                      =   1'b0;
assign   tb_i_reset[1078]                      =   1'b0;
assign   tb_i_sop[1078]                        =   1'b0;
assign   tb_i_key_update[1078]                 =   1'b0;
assign   tb_i_key[1078]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1078]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1078]               =   1'b0;
assign   tb_i_rf_static_encrypt[1078]          =   1'b1;
assign   tb_i_clear_fault_flags[1078]          =   1'b0;
assign   tb_i_rf_static_aad_length[1078]       =   64'h0000000000000100;
assign   tb_i_aad[1078]                        =   tb_i_aad[1077];
assign   tb_i_rf_static_plaintext_length[1078] =   64'h0000000000000280;
assign   tb_i_plaintext[1078]                  =   tb_i_plaintext[1077];
assign   tb_o_valid[1078]                      =   1'b0;
assign   tb_o_sop[1078]                        =   1'b0;
assign   tb_o_ciphertext[1078]                 =   tb_o_ciphertext[1077];
assign   tb_o_tag_ready[1078]                  =   1'b0;
assign   tb_o_tag[1078]                        =   tb_o_tag[1077];

// CLK no. 1079/1240
// *************************************************
assign   tb_i_valid[1079]                      =   1'b0;
assign   tb_i_reset[1079]                      =   1'b0;
assign   tb_i_sop[1079]                        =   1'b0;
assign   tb_i_key_update[1079]                 =   1'b0;
assign   tb_i_key[1079]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1079]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1079]               =   1'b0;
assign   tb_i_rf_static_encrypt[1079]          =   1'b1;
assign   tb_i_clear_fault_flags[1079]          =   1'b0;
assign   tb_i_rf_static_aad_length[1079]       =   64'h0000000000000100;
assign   tb_i_aad[1079]                        =   tb_i_aad[1078];
assign   tb_i_rf_static_plaintext_length[1079] =   64'h0000000000000280;
assign   tb_i_plaintext[1079]                  =   tb_i_plaintext[1078];
assign   tb_o_valid[1079]                      =   1'b0;
assign   tb_o_sop[1079]                        =   1'b0;
assign   tb_o_ciphertext[1079]                 =   tb_o_ciphertext[1078];
assign   tb_o_tag_ready[1079]                  =   1'b0;
assign   tb_o_tag[1079]                        =   tb_o_tag[1078];

// CLK no. 1080/1240
// *************************************************
assign   tb_i_valid[1080]                      =   1'b0;
assign   tb_i_reset[1080]                      =   1'b0;
assign   tb_i_sop[1080]                        =   1'b0;
assign   tb_i_key_update[1080]                 =   1'b0;
assign   tb_i_key[1080]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1080]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1080]               =   1'b0;
assign   tb_i_rf_static_encrypt[1080]          =   1'b1;
assign   tb_i_clear_fault_flags[1080]          =   1'b0;
assign   tb_i_rf_static_aad_length[1080]       =   64'h0000000000000100;
assign   tb_i_aad[1080]                        =   tb_i_aad[1079];
assign   tb_i_rf_static_plaintext_length[1080] =   64'h0000000000000280;
assign   tb_i_plaintext[1080]                  =   tb_i_plaintext[1079];
assign   tb_o_valid[1080]                      =   1'b0;
assign   tb_o_sop[1080]                        =   1'b0;
assign   tb_o_ciphertext[1080]                 =   tb_o_ciphertext[1079];
assign   tb_o_tag_ready[1080]                  =   1'b0;
assign   tb_o_tag[1080]                        =   tb_o_tag[1079];

// CLK no. 1081/1240
// *************************************************
assign   tb_i_valid[1081]                      =   1'b0;
assign   tb_i_reset[1081]                      =   1'b0;
assign   tb_i_sop[1081]                        =   1'b0;
assign   tb_i_key_update[1081]                 =   1'b0;
assign   tb_i_key[1081]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1081]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1081]               =   1'b0;
assign   tb_i_rf_static_encrypt[1081]          =   1'b1;
assign   tb_i_clear_fault_flags[1081]          =   1'b0;
assign   tb_i_rf_static_aad_length[1081]       =   64'h0000000000000100;
assign   tb_i_aad[1081]                        =   tb_i_aad[1080];
assign   tb_i_rf_static_plaintext_length[1081] =   64'h0000000000000280;
assign   tb_i_plaintext[1081]                  =   tb_i_plaintext[1080];
assign   tb_o_valid[1081]                      =   1'b0;
assign   tb_o_sop[1081]                        =   1'b0;
assign   tb_o_ciphertext[1081]                 =   tb_o_ciphertext[1080];
assign   tb_o_tag_ready[1081]                  =   1'b0;
assign   tb_o_tag[1081]                        =   tb_o_tag[1080];

// CLK no. 1082/1240
// *************************************************
assign   tb_i_valid[1082]                      =   1'b0;
assign   tb_i_reset[1082]                      =   1'b0;
assign   tb_i_sop[1082]                        =   1'b0;
assign   tb_i_key_update[1082]                 =   1'b0;
assign   tb_i_key[1082]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1082]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1082]               =   1'b0;
assign   tb_i_rf_static_encrypt[1082]          =   1'b1;
assign   tb_i_clear_fault_flags[1082]          =   1'b0;
assign   tb_i_rf_static_aad_length[1082]       =   64'h0000000000000100;
assign   tb_i_aad[1082]                        =   tb_i_aad[1081];
assign   tb_i_rf_static_plaintext_length[1082] =   64'h0000000000000280;
assign   tb_i_plaintext[1082]                  =   tb_i_plaintext[1081];
assign   tb_o_valid[1082]                      =   1'b0;
assign   tb_o_sop[1082]                        =   1'b0;
assign   tb_o_ciphertext[1082]                 =   tb_o_ciphertext[1081];
assign   tb_o_tag_ready[1082]                  =   1'b0;
assign   tb_o_tag[1082]                        =   tb_o_tag[1081];

// CLK no. 1083/1240
// *************************************************
assign   tb_i_valid[1083]                      =   1'b0;
assign   tb_i_reset[1083]                      =   1'b0;
assign   tb_i_sop[1083]                        =   1'b0;
assign   tb_i_key_update[1083]                 =   1'b0;
assign   tb_i_key[1083]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1083]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1083]               =   1'b0;
assign   tb_i_rf_static_encrypt[1083]          =   1'b1;
assign   tb_i_clear_fault_flags[1083]          =   1'b0;
assign   tb_i_rf_static_aad_length[1083]       =   64'h0000000000000100;
assign   tb_i_aad[1083]                        =   tb_i_aad[1082];
assign   tb_i_rf_static_plaintext_length[1083] =   64'h0000000000000280;
assign   tb_i_plaintext[1083]                  =   tb_i_plaintext[1082];
assign   tb_o_valid[1083]                      =   1'b0;
assign   tb_o_sop[1083]                        =   1'b0;
assign   tb_o_ciphertext[1083]                 =   tb_o_ciphertext[1082];
assign   tb_o_tag_ready[1083]                  =   1'b0;
assign   tb_o_tag[1083]                        =   tb_o_tag[1082];

// CLK no. 1084/1240
// *************************************************
assign   tb_i_valid[1084]                      =   1'b0;
assign   tb_i_reset[1084]                      =   1'b0;
assign   tb_i_sop[1084]                        =   1'b0;
assign   tb_i_key_update[1084]                 =   1'b0;
assign   tb_i_key[1084]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1084]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1084]               =   1'b0;
assign   tb_i_rf_static_encrypt[1084]          =   1'b1;
assign   tb_i_clear_fault_flags[1084]          =   1'b0;
assign   tb_i_rf_static_aad_length[1084]       =   64'h0000000000000100;
assign   tb_i_aad[1084]                        =   tb_i_aad[1083];
assign   tb_i_rf_static_plaintext_length[1084] =   64'h0000000000000280;
assign   tb_i_plaintext[1084]                  =   tb_i_plaintext[1083];
assign   tb_o_valid[1084]                      =   1'b0;
assign   tb_o_sop[1084]                        =   1'b0;
assign   tb_o_ciphertext[1084]                 =   tb_o_ciphertext[1083];
assign   tb_o_tag_ready[1084]                  =   1'b0;
assign   tb_o_tag[1084]                        =   tb_o_tag[1083];

// CLK no. 1085/1240
// *************************************************
assign   tb_i_valid[1085]                      =   1'b0;
assign   tb_i_reset[1085]                      =   1'b0;
assign   tb_i_sop[1085]                        =   1'b0;
assign   tb_i_key_update[1085]                 =   1'b0;
assign   tb_i_key[1085]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1085]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1085]               =   1'b0;
assign   tb_i_rf_static_encrypt[1085]          =   1'b1;
assign   tb_i_clear_fault_flags[1085]          =   1'b0;
assign   tb_i_rf_static_aad_length[1085]       =   64'h0000000000000100;
assign   tb_i_aad[1085]                        =   tb_i_aad[1084];
assign   tb_i_rf_static_plaintext_length[1085] =   64'h0000000000000280;
assign   tb_i_plaintext[1085]                  =   tb_i_plaintext[1084];
assign   tb_o_valid[1085]                      =   1'b0;
assign   tb_o_sop[1085]                        =   1'b0;
assign   tb_o_ciphertext[1085]                 =   tb_o_ciphertext[1084];
assign   tb_o_tag_ready[1085]                  =   1'b0;
assign   tb_o_tag[1085]                        =   tb_o_tag[1084];

// CLK no. 1086/1240
// *************************************************
assign   tb_i_valid[1086]                      =   1'b0;
assign   tb_i_reset[1086]                      =   1'b0;
assign   tb_i_sop[1086]                        =   1'b0;
assign   tb_i_key_update[1086]                 =   1'b0;
assign   tb_i_key[1086]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1086]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1086]               =   1'b0;
assign   tb_i_rf_static_encrypt[1086]          =   1'b1;
assign   tb_i_clear_fault_flags[1086]          =   1'b0;
assign   tb_i_rf_static_aad_length[1086]       =   64'h0000000000000100;
assign   tb_i_aad[1086]                        =   tb_i_aad[1085];
assign   tb_i_rf_static_plaintext_length[1086] =   64'h0000000000000280;
assign   tb_i_plaintext[1086]                  =   tb_i_plaintext[1085];
assign   tb_o_valid[1086]                      =   1'b0;
assign   tb_o_sop[1086]                        =   1'b0;
assign   tb_o_ciphertext[1086]                 =   tb_o_ciphertext[1085];
assign   tb_o_tag_ready[1086]                  =   1'b0;
assign   tb_o_tag[1086]                        =   tb_o_tag[1085];

// CLK no. 1087/1240
// *************************************************
assign   tb_i_valid[1087]                      =   1'b0;
assign   tb_i_reset[1087]                      =   1'b0;
assign   tb_i_sop[1087]                        =   1'b0;
assign   tb_i_key_update[1087]                 =   1'b0;
assign   tb_i_key[1087]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1087]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1087]               =   1'b0;
assign   tb_i_rf_static_encrypt[1087]          =   1'b1;
assign   tb_i_clear_fault_flags[1087]          =   1'b0;
assign   tb_i_rf_static_aad_length[1087]       =   64'h0000000000000100;
assign   tb_i_aad[1087]                        =   tb_i_aad[1086];
assign   tb_i_rf_static_plaintext_length[1087] =   64'h0000000000000280;
assign   tb_i_plaintext[1087]                  =   tb_i_plaintext[1086];
assign   tb_o_valid[1087]                      =   1'b0;
assign   tb_o_sop[1087]                        =   1'b0;
assign   tb_o_ciphertext[1087]                 =   tb_o_ciphertext[1086];
assign   tb_o_tag_ready[1087]                  =   1'b0;
assign   tb_o_tag[1087]                        =   tb_o_tag[1086];

// CLK no. 1088/1240
// *************************************************
assign   tb_i_valid[1088]                      =   1'b0;
assign   tb_i_reset[1088]                      =   1'b0;
assign   tb_i_sop[1088]                        =   1'b0;
assign   tb_i_key_update[1088]                 =   1'b0;
assign   tb_i_key[1088]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1088]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1088]               =   1'b0;
assign   tb_i_rf_static_encrypt[1088]          =   1'b1;
assign   tb_i_clear_fault_flags[1088]          =   1'b0;
assign   tb_i_rf_static_aad_length[1088]       =   64'h0000000000000100;
assign   tb_i_aad[1088]                        =   tb_i_aad[1087];
assign   tb_i_rf_static_plaintext_length[1088] =   64'h0000000000000280;
assign   tb_i_plaintext[1088]                  =   tb_i_plaintext[1087];
assign   tb_o_valid[1088]                      =   1'b0;
assign   tb_o_sop[1088]                        =   1'b0;
assign   tb_o_ciphertext[1088]                 =   tb_o_ciphertext[1087];
assign   tb_o_tag_ready[1088]                  =   1'b0;
assign   tb_o_tag[1088]                        =   tb_o_tag[1087];

// CLK no. 1089/1240
// *************************************************
assign   tb_i_valid[1089]                      =   1'b0;
assign   tb_i_reset[1089]                      =   1'b0;
assign   tb_i_sop[1089]                        =   1'b0;
assign   tb_i_key_update[1089]                 =   1'b0;
assign   tb_i_key[1089]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1089]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1089]               =   1'b0;
assign   tb_i_rf_static_encrypt[1089]          =   1'b1;
assign   tb_i_clear_fault_flags[1089]          =   1'b0;
assign   tb_i_rf_static_aad_length[1089]       =   64'h0000000000000100;
assign   tb_i_aad[1089]                        =   tb_i_aad[1088];
assign   tb_i_rf_static_plaintext_length[1089] =   64'h0000000000000280;
assign   tb_i_plaintext[1089]                  =   tb_i_plaintext[1088];
assign   tb_o_valid[1089]                      =   1'b0;
assign   tb_o_sop[1089]                        =   1'b0;
assign   tb_o_ciphertext[1089]                 =   tb_o_ciphertext[1088];
assign   tb_o_tag_ready[1089]                  =   1'b0;
assign   tb_o_tag[1089]                        =   tb_o_tag[1088];

// CLK no. 1090/1240
// *************************************************
assign   tb_i_valid[1090]                      =   1'b0;
assign   tb_i_reset[1090]                      =   1'b0;
assign   tb_i_sop[1090]                        =   1'b0;
assign   tb_i_key_update[1090]                 =   1'b0;
assign   tb_i_key[1090]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1090]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1090]               =   1'b0;
assign   tb_i_rf_static_encrypt[1090]          =   1'b1;
assign   tb_i_clear_fault_flags[1090]          =   1'b0;
assign   tb_i_rf_static_aad_length[1090]       =   64'h0000000000000100;
assign   tb_i_aad[1090]                        =   tb_i_aad[1089];
assign   tb_i_rf_static_plaintext_length[1090] =   64'h0000000000000280;
assign   tb_i_plaintext[1090]                  =   tb_i_plaintext[1089];
assign   tb_o_valid[1090]                      =   1'b0;
assign   tb_o_sop[1090]                        =   1'b0;
assign   tb_o_ciphertext[1090]                 =   tb_o_ciphertext[1089];
assign   tb_o_tag_ready[1090]                  =   1'b0;
assign   tb_o_tag[1090]                        =   tb_o_tag[1089];

// CLK no. 1091/1240
// *************************************************
assign   tb_i_valid[1091]                      =   1'b0;
assign   tb_i_reset[1091]                      =   1'b0;
assign   tb_i_sop[1091]                        =   1'b0;
assign   tb_i_key_update[1091]                 =   1'b0;
assign   tb_i_key[1091]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1091]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1091]               =   1'b0;
assign   tb_i_rf_static_encrypt[1091]          =   1'b1;
assign   tb_i_clear_fault_flags[1091]          =   1'b0;
assign   tb_i_rf_static_aad_length[1091]       =   64'h0000000000000100;
assign   tb_i_aad[1091]                        =   tb_i_aad[1090];
assign   tb_i_rf_static_plaintext_length[1091] =   64'h0000000000000280;
assign   tb_i_plaintext[1091]                  =   tb_i_plaintext[1090];
assign   tb_o_valid[1091]                      =   1'b0;
assign   tb_o_sop[1091]                        =   1'b0;
assign   tb_o_ciphertext[1091]                 =   tb_o_ciphertext[1090];
assign   tb_o_tag_ready[1091]                  =   1'b0;
assign   tb_o_tag[1091]                        =   tb_o_tag[1090];

// CLK no. 1092/1240
// *************************************************
assign   tb_i_valid[1092]                      =   1'b0;
assign   tb_i_reset[1092]                      =   1'b0;
assign   tb_i_sop[1092]                        =   1'b0;
assign   tb_i_key_update[1092]                 =   1'b0;
assign   tb_i_key[1092]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1092]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1092]               =   1'b0;
assign   tb_i_rf_static_encrypt[1092]          =   1'b1;
assign   tb_i_clear_fault_flags[1092]          =   1'b0;
assign   tb_i_rf_static_aad_length[1092]       =   64'h0000000000000100;
assign   tb_i_aad[1092]                        =   tb_i_aad[1091];
assign   tb_i_rf_static_plaintext_length[1092] =   64'h0000000000000280;
assign   tb_i_plaintext[1092]                  =   tb_i_plaintext[1091];
assign   tb_o_valid[1092]                      =   1'b0;
assign   tb_o_sop[1092]                        =   1'b0;
assign   tb_o_ciphertext[1092]                 =   tb_o_ciphertext[1091];
assign   tb_o_tag_ready[1092]                  =   1'b0;
assign   tb_o_tag[1092]                        =   tb_o_tag[1091];

// CLK no. 1093/1240
// *************************************************
assign   tb_i_valid[1093]                      =   1'b0;
assign   tb_i_reset[1093]                      =   1'b0;
assign   tb_i_sop[1093]                        =   1'b0;
assign   tb_i_key_update[1093]                 =   1'b0;
assign   tb_i_key[1093]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1093]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1093]               =   1'b0;
assign   tb_i_rf_static_encrypt[1093]          =   1'b1;
assign   tb_i_clear_fault_flags[1093]          =   1'b0;
assign   tb_i_rf_static_aad_length[1093]       =   64'h0000000000000100;
assign   tb_i_aad[1093]                        =   tb_i_aad[1092];
assign   tb_i_rf_static_plaintext_length[1093] =   64'h0000000000000280;
assign   tb_i_plaintext[1093]                  =   tb_i_plaintext[1092];
assign   tb_o_valid[1093]                      =   1'b0;
assign   tb_o_sop[1093]                        =   1'b0;
assign   tb_o_ciphertext[1093]                 =   tb_o_ciphertext[1092];
assign   tb_o_tag_ready[1093]                  =   1'b0;
assign   tb_o_tag[1093]                        =   tb_o_tag[1092];

// CLK no. 1094/1240
// *************************************************
assign   tb_i_valid[1094]                      =   1'b0;
assign   tb_i_reset[1094]                      =   1'b0;
assign   tb_i_sop[1094]                        =   1'b0;
assign   tb_i_key_update[1094]                 =   1'b0;
assign   tb_i_key[1094]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1094]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1094]               =   1'b0;
assign   tb_i_rf_static_encrypt[1094]          =   1'b1;
assign   tb_i_clear_fault_flags[1094]          =   1'b0;
assign   tb_i_rf_static_aad_length[1094]       =   64'h0000000000000100;
assign   tb_i_aad[1094]                        =   tb_i_aad[1093];
assign   tb_i_rf_static_plaintext_length[1094] =   64'h0000000000000280;
assign   tb_i_plaintext[1094]                  =   tb_i_plaintext[1093];
assign   tb_o_valid[1094]                      =   1'b0;
assign   tb_o_sop[1094]                        =   1'b0;
assign   tb_o_ciphertext[1094]                 =   tb_o_ciphertext[1093];
assign   tb_o_tag_ready[1094]                  =   1'b0;
assign   tb_o_tag[1094]                        =   tb_o_tag[1093];

// CLK no. 1095/1240
// *************************************************
assign   tb_i_valid[1095]                      =   1'b0;
assign   tb_i_reset[1095]                      =   1'b0;
assign   tb_i_sop[1095]                        =   1'b0;
assign   tb_i_key_update[1095]                 =   1'b0;
assign   tb_i_key[1095]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1095]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1095]               =   1'b0;
assign   tb_i_rf_static_encrypt[1095]          =   1'b1;
assign   tb_i_clear_fault_flags[1095]          =   1'b0;
assign   tb_i_rf_static_aad_length[1095]       =   64'h0000000000000100;
assign   tb_i_aad[1095]                        =   tb_i_aad[1094];
assign   tb_i_rf_static_plaintext_length[1095] =   64'h0000000000000280;
assign   tb_i_plaintext[1095]                  =   tb_i_plaintext[1094];
assign   tb_o_valid[1095]                      =   1'b0;
assign   tb_o_sop[1095]                        =   1'b0;
assign   tb_o_ciphertext[1095]                 =   tb_o_ciphertext[1094];
assign   tb_o_tag_ready[1095]                  =   1'b0;
assign   tb_o_tag[1095]                        =   tb_o_tag[1094];

// CLK no. 1096/1240
// *************************************************
assign   tb_i_valid[1096]                      =   1'b0;
assign   tb_i_reset[1096]                      =   1'b0;
assign   tb_i_sop[1096]                        =   1'b0;
assign   tb_i_key_update[1096]                 =   1'b0;
assign   tb_i_key[1096]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1096]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1096]               =   1'b0;
assign   tb_i_rf_static_encrypt[1096]          =   1'b1;
assign   tb_i_clear_fault_flags[1096]          =   1'b0;
assign   tb_i_rf_static_aad_length[1096]       =   64'h0000000000000100;
assign   tb_i_aad[1096]                        =   tb_i_aad[1095];
assign   tb_i_rf_static_plaintext_length[1096] =   64'h0000000000000280;
assign   tb_i_plaintext[1096]                  =   tb_i_plaintext[1095];
assign   tb_o_valid[1096]                      =   1'b0;
assign   tb_o_sop[1096]                        =   1'b0;
assign   tb_o_ciphertext[1096]                 =   tb_o_ciphertext[1095];
assign   tb_o_tag_ready[1096]                  =   1'b0;
assign   tb_o_tag[1096]                        =   tb_o_tag[1095];

// CLK no. 1097/1240
// *************************************************
assign   tb_i_valid[1097]                      =   1'b0;
assign   tb_i_reset[1097]                      =   1'b0;
assign   tb_i_sop[1097]                        =   1'b0;
assign   tb_i_key_update[1097]                 =   1'b0;
assign   tb_i_key[1097]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1097]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1097]               =   1'b0;
assign   tb_i_rf_static_encrypt[1097]          =   1'b1;
assign   tb_i_clear_fault_flags[1097]          =   1'b0;
assign   tb_i_rf_static_aad_length[1097]       =   64'h0000000000000100;
assign   tb_i_aad[1097]                        =   tb_i_aad[1096];
assign   tb_i_rf_static_plaintext_length[1097] =   64'h0000000000000280;
assign   tb_i_plaintext[1097]                  =   tb_i_plaintext[1096];
assign   tb_o_valid[1097]                      =   1'b0;
assign   tb_o_sop[1097]                        =   1'b0;
assign   tb_o_ciphertext[1097]                 =   tb_o_ciphertext[1096];
assign   tb_o_tag_ready[1097]                  =   1'b0;
assign   tb_o_tag[1097]                        =   tb_o_tag[1096];

// CLK no. 1098/1240
// *************************************************
assign   tb_i_valid[1098]                      =   1'b0;
assign   tb_i_reset[1098]                      =   1'b0;
assign   tb_i_sop[1098]                        =   1'b0;
assign   tb_i_key_update[1098]                 =   1'b0;
assign   tb_i_key[1098]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1098]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1098]               =   1'b0;
assign   tb_i_rf_static_encrypt[1098]          =   1'b1;
assign   tb_i_clear_fault_flags[1098]          =   1'b0;
assign   tb_i_rf_static_aad_length[1098]       =   64'h0000000000000100;
assign   tb_i_aad[1098]                        =   tb_i_aad[1097];
assign   tb_i_rf_static_plaintext_length[1098] =   64'h0000000000000280;
assign   tb_i_plaintext[1098]                  =   tb_i_plaintext[1097];
assign   tb_o_valid[1098]                      =   1'b0;
assign   tb_o_sop[1098]                        =   1'b0;
assign   tb_o_ciphertext[1098]                 =   tb_o_ciphertext[1097];
assign   tb_o_tag_ready[1098]                  =   1'b0;
assign   tb_o_tag[1098]                        =   tb_o_tag[1097];

// CLK no. 1099/1240
// *************************************************
assign   tb_i_valid[1099]                      =   1'b0;
assign   tb_i_reset[1099]                      =   1'b0;
assign   tb_i_sop[1099]                        =   1'b0;
assign   tb_i_key_update[1099]                 =   1'b0;
assign   tb_i_key[1099]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1099]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1099]               =   1'b0;
assign   tb_i_rf_static_encrypt[1099]          =   1'b1;
assign   tb_i_clear_fault_flags[1099]          =   1'b0;
assign   tb_i_rf_static_aad_length[1099]       =   64'h0000000000000100;
assign   tb_i_aad[1099]                        =   tb_i_aad[1098];
assign   tb_i_rf_static_plaintext_length[1099] =   64'h0000000000000280;
assign   tb_i_plaintext[1099]                  =   tb_i_plaintext[1098];
assign   tb_o_valid[1099]                      =   1'b0;
assign   tb_o_sop[1099]                        =   1'b0;
assign   tb_o_ciphertext[1099]                 =   tb_o_ciphertext[1098];
assign   tb_o_tag_ready[1099]                  =   1'b0;
assign   tb_o_tag[1099]                        =   tb_o_tag[1098];

// CLK no. 1100/1240
// *************************************************
assign   tb_i_valid[1100]                      =   1'b0;
assign   tb_i_reset[1100]                      =   1'b0;
assign   tb_i_sop[1100]                        =   1'b0;
assign   tb_i_key_update[1100]                 =   1'b0;
assign   tb_i_key[1100]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1100]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1100]               =   1'b0;
assign   tb_i_rf_static_encrypt[1100]          =   1'b1;
assign   tb_i_clear_fault_flags[1100]          =   1'b0;
assign   tb_i_rf_static_aad_length[1100]       =   64'h0000000000000100;
assign   tb_i_aad[1100]                        =   tb_i_aad[1099];
assign   tb_i_rf_static_plaintext_length[1100] =   64'h0000000000000280;
assign   tb_i_plaintext[1100]                  =   tb_i_plaintext[1099];
assign   tb_o_valid[1100]                      =   1'b0;
assign   tb_o_sop[1100]                        =   1'b0;
assign   tb_o_ciphertext[1100]                 =   tb_o_ciphertext[1099];
assign   tb_o_tag_ready[1100]                  =   1'b0;
assign   tb_o_tag[1100]                        =   tb_o_tag[1099];

// CLK no. 1101/1240
// *************************************************
assign   tb_i_valid[1101]                      =   1'b0;
assign   tb_i_reset[1101]                      =   1'b0;
assign   tb_i_sop[1101]                        =   1'b0;
assign   tb_i_key_update[1101]                 =   1'b0;
assign   tb_i_key[1101]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1101]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1101]               =   1'b0;
assign   tb_i_rf_static_encrypt[1101]          =   1'b1;
assign   tb_i_clear_fault_flags[1101]          =   1'b0;
assign   tb_i_rf_static_aad_length[1101]       =   64'h0000000000000100;
assign   tb_i_aad[1101]                        =   tb_i_aad[1100];
assign   tb_i_rf_static_plaintext_length[1101] =   64'h0000000000000280;
assign   tb_i_plaintext[1101]                  =   tb_i_plaintext[1100];
assign   tb_o_valid[1101]                      =   1'b0;
assign   tb_o_sop[1101]                        =   1'b0;
assign   tb_o_ciphertext[1101]                 =   tb_o_ciphertext[1100];
assign   tb_o_tag_ready[1101]                  =   1'b0;
assign   tb_o_tag[1101]                        =   tb_o_tag[1100];

// CLK no. 1102/1240
// *************************************************
assign   tb_i_valid[1102]                      =   1'b0;
assign   tb_i_reset[1102]                      =   1'b0;
assign   tb_i_sop[1102]                        =   1'b0;
assign   tb_i_key_update[1102]                 =   1'b0;
assign   tb_i_key[1102]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1102]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1102]               =   1'b0;
assign   tb_i_rf_static_encrypt[1102]          =   1'b1;
assign   tb_i_clear_fault_flags[1102]          =   1'b0;
assign   tb_i_rf_static_aad_length[1102]       =   64'h0000000000000100;
assign   tb_i_aad[1102]                        =   tb_i_aad[1101];
assign   tb_i_rf_static_plaintext_length[1102] =   64'h0000000000000280;
assign   tb_i_plaintext[1102]                  =   tb_i_plaintext[1101];
assign   tb_o_valid[1102]                      =   1'b0;
assign   tb_o_sop[1102]                        =   1'b0;
assign   tb_o_ciphertext[1102]                 =   tb_o_ciphertext[1101];
assign   tb_o_tag_ready[1102]                  =   1'b0;
assign   tb_o_tag[1102]                        =   tb_o_tag[1101];

// CLK no. 1103/1240
// *************************************************
assign   tb_i_valid[1103]                      =   1'b0;
assign   tb_i_reset[1103]                      =   1'b0;
assign   tb_i_sop[1103]                        =   1'b0;
assign   tb_i_key_update[1103]                 =   1'b0;
assign   tb_i_key[1103]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1103]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1103]               =   1'b0;
assign   tb_i_rf_static_encrypt[1103]          =   1'b1;
assign   tb_i_clear_fault_flags[1103]          =   1'b0;
assign   tb_i_rf_static_aad_length[1103]       =   64'h0000000000000100;
assign   tb_i_aad[1103]                        =   tb_i_aad[1102];
assign   tb_i_rf_static_plaintext_length[1103] =   64'h0000000000000280;
assign   tb_i_plaintext[1103]                  =   tb_i_plaintext[1102];
assign   tb_o_valid[1103]                      =   1'b0;
assign   tb_o_sop[1103]                        =   1'b0;
assign   tb_o_ciphertext[1103]                 =   tb_o_ciphertext[1102];
assign   tb_o_tag_ready[1103]                  =   1'b0;
assign   tb_o_tag[1103]                        =   tb_o_tag[1102];

// CLK no. 1104/1240
// *************************************************
assign   tb_i_valid[1104]                      =   1'b0;
assign   tb_i_reset[1104]                      =   1'b0;
assign   tb_i_sop[1104]                        =   1'b0;
assign   tb_i_key_update[1104]                 =   1'b0;
assign   tb_i_key[1104]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1104]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1104]               =   1'b0;
assign   tb_i_rf_static_encrypt[1104]          =   1'b1;
assign   tb_i_clear_fault_flags[1104]          =   1'b0;
assign   tb_i_rf_static_aad_length[1104]       =   64'h0000000000000100;
assign   tb_i_aad[1104]                        =   tb_i_aad[1103];
assign   tb_i_rf_static_plaintext_length[1104] =   64'h0000000000000280;
assign   tb_i_plaintext[1104]                  =   tb_i_plaintext[1103];
assign   tb_o_valid[1104]                      =   1'b0;
assign   tb_o_sop[1104]                        =   1'b0;
assign   tb_o_ciphertext[1104]                 =   tb_o_ciphertext[1103];
assign   tb_o_tag_ready[1104]                  =   1'b0;
assign   tb_o_tag[1104]                        =   tb_o_tag[1103];

// CLK no. 1105/1240
// *************************************************
assign   tb_i_valid[1105]                      =   1'b0;
assign   tb_i_reset[1105]                      =   1'b0;
assign   tb_i_sop[1105]                        =   1'b0;
assign   tb_i_key_update[1105]                 =   1'b0;
assign   tb_i_key[1105]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1105]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1105]               =   1'b0;
assign   tb_i_rf_static_encrypt[1105]          =   1'b1;
assign   tb_i_clear_fault_flags[1105]          =   1'b0;
assign   tb_i_rf_static_aad_length[1105]       =   64'h0000000000000100;
assign   tb_i_aad[1105]                        =   tb_i_aad[1104];
assign   tb_i_rf_static_plaintext_length[1105] =   64'h0000000000000280;
assign   tb_i_plaintext[1105]                  =   tb_i_plaintext[1104];
assign   tb_o_valid[1105]                      =   1'b0;
assign   tb_o_sop[1105]                        =   1'b0;
assign   tb_o_ciphertext[1105]                 =   tb_o_ciphertext[1104];
assign   tb_o_tag_ready[1105]                  =   1'b0;
assign   tb_o_tag[1105]                        =   tb_o_tag[1104];

// CLK no. 1106/1240
// *************************************************
assign   tb_i_valid[1106]                      =   1'b0;
assign   tb_i_reset[1106]                      =   1'b0;
assign   tb_i_sop[1106]                        =   1'b0;
assign   tb_i_key_update[1106]                 =   1'b0;
assign   tb_i_key[1106]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1106]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1106]               =   1'b0;
assign   tb_i_rf_static_encrypt[1106]          =   1'b1;
assign   tb_i_clear_fault_flags[1106]          =   1'b0;
assign   tb_i_rf_static_aad_length[1106]       =   64'h0000000000000100;
assign   tb_i_aad[1106]                        =   tb_i_aad[1105];
assign   tb_i_rf_static_plaintext_length[1106] =   64'h0000000000000280;
assign   tb_i_plaintext[1106]                  =   tb_i_plaintext[1105];
assign   tb_o_valid[1106]                      =   1'b0;
assign   tb_o_sop[1106]                        =   1'b0;
assign   tb_o_ciphertext[1106]                 =   tb_o_ciphertext[1105];
assign   tb_o_tag_ready[1106]                  =   1'b0;
assign   tb_o_tag[1106]                        =   tb_o_tag[1105];

// CLK no. 1107/1240
// *************************************************
assign   tb_i_valid[1107]                      =   1'b0;
assign   tb_i_reset[1107]                      =   1'b0;
assign   tb_i_sop[1107]                        =   1'b0;
assign   tb_i_key_update[1107]                 =   1'b0;
assign   tb_i_key[1107]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1107]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1107]               =   1'b0;
assign   tb_i_rf_static_encrypt[1107]          =   1'b1;
assign   tb_i_clear_fault_flags[1107]          =   1'b0;
assign   tb_i_rf_static_aad_length[1107]       =   64'h0000000000000100;
assign   tb_i_aad[1107]                        =   tb_i_aad[1106];
assign   tb_i_rf_static_plaintext_length[1107] =   64'h0000000000000280;
assign   tb_i_plaintext[1107]                  =   tb_i_plaintext[1106];
assign   tb_o_valid[1107]                      =   1'b0;
assign   tb_o_sop[1107]                        =   1'b0;
assign   tb_o_ciphertext[1107]                 =   tb_o_ciphertext[1106];
assign   tb_o_tag_ready[1107]                  =   1'b0;
assign   tb_o_tag[1107]                        =   tb_o_tag[1106];

// CLK no. 1108/1240
// *************************************************
assign   tb_i_valid[1108]                      =   1'b0;
assign   tb_i_reset[1108]                      =   1'b0;
assign   tb_i_sop[1108]                        =   1'b0;
assign   tb_i_key_update[1108]                 =   1'b0;
assign   tb_i_key[1108]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1108]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1108]               =   1'b0;
assign   tb_i_rf_static_encrypt[1108]          =   1'b1;
assign   tb_i_clear_fault_flags[1108]          =   1'b0;
assign   tb_i_rf_static_aad_length[1108]       =   64'h0000000000000100;
assign   tb_i_aad[1108]                        =   tb_i_aad[1107];
assign   tb_i_rf_static_plaintext_length[1108] =   64'h0000000000000280;
assign   tb_i_plaintext[1108]                  =   tb_i_plaintext[1107];
assign   tb_o_valid[1108]                      =   1'b0;
assign   tb_o_sop[1108]                        =   1'b0;
assign   tb_o_ciphertext[1108]                 =   tb_o_ciphertext[1107];
assign   tb_o_tag_ready[1108]                  =   1'b0;
assign   tb_o_tag[1108]                        =   tb_o_tag[1107];

// CLK no. 1109/1240
// *************************************************
assign   tb_i_valid[1109]                      =   1'b0;
assign   tb_i_reset[1109]                      =   1'b0;
assign   tb_i_sop[1109]                        =   1'b0;
assign   tb_i_key_update[1109]                 =   1'b0;
assign   tb_i_key[1109]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1109]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1109]               =   1'b0;
assign   tb_i_rf_static_encrypt[1109]          =   1'b1;
assign   tb_i_clear_fault_flags[1109]          =   1'b0;
assign   tb_i_rf_static_aad_length[1109]       =   64'h0000000000000100;
assign   tb_i_aad[1109]                        =   tb_i_aad[1108];
assign   tb_i_rf_static_plaintext_length[1109] =   64'h0000000000000280;
assign   tb_i_plaintext[1109]                  =   tb_i_plaintext[1108];
assign   tb_o_valid[1109]                      =   1'b1;
assign   tb_o_sop[1109]                        =   1'b1;
assign   tb_o_ciphertext[1109]                 =   256'h191866921edfca4cf58916c64b21d597be33e4d2b4493cba961c11c8c5108003;
assign   tb_o_tag_ready[1109]                  =   1'b0;
assign   tb_o_tag[1109]                        =   tb_o_tag[1108];

// CLK no. 1110/1240
// *************************************************
assign   tb_i_valid[1110]                      =   1'b0;
assign   tb_i_reset[1110]                      =   1'b0;
assign   tb_i_sop[1110]                        =   1'b0;
assign   tb_i_key_update[1110]                 =   1'b0;
assign   tb_i_key[1110]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1110]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1110]               =   1'b0;
assign   tb_i_rf_static_encrypt[1110]          =   1'b1;
assign   tb_i_clear_fault_flags[1110]          =   1'b0;
assign   tb_i_rf_static_aad_length[1110]       =   64'h0000000000000100;
assign   tb_i_aad[1110]                        =   tb_i_aad[1109];
assign   tb_i_rf_static_plaintext_length[1110] =   64'h0000000000000280;
assign   tb_i_plaintext[1110]                  =   tb_i_plaintext[1109];
assign   tb_o_valid[1110]                      =   1'b1;
assign   tb_o_sop[1110]                        =   1'b0;
assign   tb_o_ciphertext[1110]                 =   256'h06fd7fa9eeff6fa5af0a40021925b81f9910bf2ddac4e65861a9cff1abc0c07d;
assign   tb_o_tag_ready[1110]                  =   1'b0;
assign   tb_o_tag[1110]                        =   tb_o_tag[1109];

// CLK no. 1111/1240
// *************************************************
assign   tb_i_valid[1111]                      =   1'b0;
assign   tb_i_reset[1111]                      =   1'b0;
assign   tb_i_sop[1111]                        =   1'b0;
assign   tb_i_key_update[1111]                 =   1'b0;
assign   tb_i_key[1111]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1111]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1111]               =   1'b0;
assign   tb_i_rf_static_encrypt[1111]          =   1'b1;
assign   tb_i_clear_fault_flags[1111]          =   1'b0;
assign   tb_i_rf_static_aad_length[1111]       =   64'h0000000000000100;
assign   tb_i_aad[1111]                        =   tb_i_aad[1110];
assign   tb_i_rf_static_plaintext_length[1111] =   64'h0000000000000280;
assign   tb_i_plaintext[1111]                  =   tb_i_plaintext[1110];
assign   tb_o_valid[1111]                      =   1'b1;
assign   tb_o_sop[1111]                        =   1'b0;
assign   tb_o_ciphertext[1111]                 =   256'h91456498128b0ddeca448d8cb8f61f2d;
assign   tb_o_tag_ready[1111]                  =   1'b0;
assign   tb_o_tag[1111]                        =   tb_o_tag[1110];

// CLK no. 1112/1240
// *************************************************
assign   tb_i_valid[1112]                      =   1'b0;
assign   tb_i_reset[1112]                      =   1'b0;
assign   tb_i_sop[1112]                        =   1'b0;
assign   tb_i_key_update[1112]                 =   1'b0;
assign   tb_i_key[1112]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1112]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1112]               =   1'b0;
assign   tb_i_rf_static_encrypt[1112]          =   1'b1;
assign   tb_i_clear_fault_flags[1112]          =   1'b0;
assign   tb_i_rf_static_aad_length[1112]       =   64'h0000000000000100;
assign   tb_i_aad[1112]                        =   tb_i_aad[1111];
assign   tb_i_rf_static_plaintext_length[1112] =   64'h0000000000000280;
assign   tb_i_plaintext[1112]                  =   tb_i_plaintext[1111];
assign   tb_o_valid[1112]                      =   1'b0;
assign   tb_o_sop[1112]                        =   1'b0;
assign   tb_o_ciphertext[1112]                 =   tb_o_ciphertext[1111];
assign   tb_o_tag_ready[1112]                  =   1'b0;
assign   tb_o_tag[1112]                        =   tb_o_tag[1111];

// CLK no. 1113/1240
// *************************************************
assign   tb_i_valid[1113]                      =   1'b0;
assign   tb_i_reset[1113]                      =   1'b0;
assign   tb_i_sop[1113]                        =   1'b0;
assign   tb_i_key_update[1113]                 =   1'b0;
assign   tb_i_key[1113]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1113]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1113]               =   1'b0;
assign   tb_i_rf_static_encrypt[1113]          =   1'b1;
assign   tb_i_clear_fault_flags[1113]          =   1'b0;
assign   tb_i_rf_static_aad_length[1113]       =   64'h0000000000000100;
assign   tb_i_aad[1113]                        =   tb_i_aad[1112];
assign   tb_i_rf_static_plaintext_length[1113] =   64'h0000000000000280;
assign   tb_i_plaintext[1113]                  =   tb_i_plaintext[1112];
assign   tb_o_valid[1113]                      =   1'b0;
assign   tb_o_sop[1113]                        =   1'b0;
assign   tb_o_ciphertext[1113]                 =   tb_o_ciphertext[1112];
assign   tb_o_tag_ready[1113]                  =   1'b0;
assign   tb_o_tag[1113]                        =   tb_o_tag[1112];

// CLK no. 1114/1240
// *************************************************
assign   tb_i_valid[1114]                      =   1'b0;
assign   tb_i_reset[1114]                      =   1'b0;
assign   tb_i_sop[1114]                        =   1'b0;
assign   tb_i_key_update[1114]                 =   1'b0;
assign   tb_i_key[1114]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1114]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1114]               =   1'b0;
assign   tb_i_rf_static_encrypt[1114]          =   1'b1;
assign   tb_i_clear_fault_flags[1114]          =   1'b0;
assign   tb_i_rf_static_aad_length[1114]       =   64'h0000000000000100;
assign   tb_i_aad[1114]                        =   tb_i_aad[1113];
assign   tb_i_rf_static_plaintext_length[1114] =   64'h0000000000000280;
assign   tb_i_plaintext[1114]                  =   tb_i_plaintext[1113];
assign   tb_o_valid[1114]                      =   1'b0;
assign   tb_o_sop[1114]                        =   1'b0;
assign   tb_o_ciphertext[1114]                 =   tb_o_ciphertext[1113];
assign   tb_o_tag_ready[1114]                  =   1'b0;
assign   tb_o_tag[1114]                        =   tb_o_tag[1113];

// CLK no. 1115/1240
// *************************************************
assign   tb_i_valid[1115]                      =   1'b0;
assign   tb_i_reset[1115]                      =   1'b0;
assign   tb_i_sop[1115]                        =   1'b0;
assign   tb_i_key_update[1115]                 =   1'b0;
assign   tb_i_key[1115]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1115]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1115]               =   1'b0;
assign   tb_i_rf_static_encrypt[1115]          =   1'b1;
assign   tb_i_clear_fault_flags[1115]          =   1'b0;
assign   tb_i_rf_static_aad_length[1115]       =   64'h0000000000000100;
assign   tb_i_aad[1115]                        =   tb_i_aad[1114];
assign   tb_i_rf_static_plaintext_length[1115] =   64'h0000000000000280;
assign   tb_i_plaintext[1115]                  =   tb_i_plaintext[1114];
assign   tb_o_valid[1115]                      =   1'b0;
assign   tb_o_sop[1115]                        =   1'b0;
assign   tb_o_ciphertext[1115]                 =   tb_o_ciphertext[1114];
assign   tb_o_tag_ready[1115]                  =   1'b0;
assign   tb_o_tag[1115]                        =   tb_o_tag[1114];

// CLK no. 1116/1240
// *************************************************
assign   tb_i_valid[1116]                      =   1'b0;
assign   tb_i_reset[1116]                      =   1'b0;
assign   tb_i_sop[1116]                        =   1'b0;
assign   tb_i_key_update[1116]                 =   1'b0;
assign   tb_i_key[1116]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1116]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1116]               =   1'b0;
assign   tb_i_rf_static_encrypt[1116]          =   1'b1;
assign   tb_i_clear_fault_flags[1116]          =   1'b0;
assign   tb_i_rf_static_aad_length[1116]       =   64'h0000000000000100;
assign   tb_i_aad[1116]                        =   tb_i_aad[1115];
assign   tb_i_rf_static_plaintext_length[1116] =   64'h0000000000000280;
assign   tb_i_plaintext[1116]                  =   tb_i_plaintext[1115];
assign   tb_o_valid[1116]                      =   1'b0;
assign   tb_o_sop[1116]                        =   1'b0;
assign   tb_o_ciphertext[1116]                 =   tb_o_ciphertext[1115];
assign   tb_o_tag_ready[1116]                  =   1'b0;
assign   tb_o_tag[1116]                        =   tb_o_tag[1115];

// CLK no. 1117/1240
// *************************************************
assign   tb_i_valid[1117]                      =   1'b0;
assign   tb_i_reset[1117]                      =   1'b0;
assign   tb_i_sop[1117]                        =   1'b0;
assign   tb_i_key_update[1117]                 =   1'b0;
assign   tb_i_key[1117]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1117]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1117]               =   1'b0;
assign   tb_i_rf_static_encrypt[1117]          =   1'b1;
assign   tb_i_clear_fault_flags[1117]          =   1'b0;
assign   tb_i_rf_static_aad_length[1117]       =   64'h0000000000000100;
assign   tb_i_aad[1117]                        =   tb_i_aad[1116];
assign   tb_i_rf_static_plaintext_length[1117] =   64'h0000000000000280;
assign   tb_i_plaintext[1117]                  =   tb_i_plaintext[1116];
assign   tb_o_valid[1117]                      =   1'b0;
assign   tb_o_sop[1117]                        =   1'b0;
assign   tb_o_ciphertext[1117]                 =   tb_o_ciphertext[1116];
assign   tb_o_tag_ready[1117]                  =   1'b0;
assign   tb_o_tag[1117]                        =   tb_o_tag[1116];

// CLK no. 1118/1240
// *************************************************
assign   tb_i_valid[1118]                      =   1'b0;
assign   tb_i_reset[1118]                      =   1'b0;
assign   tb_i_sop[1118]                        =   1'b0;
assign   tb_i_key_update[1118]                 =   1'b0;
assign   tb_i_key[1118]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1118]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1118]               =   1'b0;
assign   tb_i_rf_static_encrypt[1118]          =   1'b1;
assign   tb_i_clear_fault_flags[1118]          =   1'b0;
assign   tb_i_rf_static_aad_length[1118]       =   64'h0000000000000100;
assign   tb_i_aad[1118]                        =   tb_i_aad[1117];
assign   tb_i_rf_static_plaintext_length[1118] =   64'h0000000000000280;
assign   tb_i_plaintext[1118]                  =   tb_i_plaintext[1117];
assign   tb_o_valid[1118]                      =   1'b0;
assign   tb_o_sop[1118]                        =   1'b0;
assign   tb_o_ciphertext[1118]                 =   tb_o_ciphertext[1117];
assign   tb_o_tag_ready[1118]                  =   1'b0;
assign   tb_o_tag[1118]                        =   tb_o_tag[1117];

// CLK no. 1119/1240
// *************************************************
assign   tb_i_valid[1119]                      =   1'b0;
assign   tb_i_reset[1119]                      =   1'b0;
assign   tb_i_sop[1119]                        =   1'b0;
assign   tb_i_key_update[1119]                 =   1'b0;
assign   tb_i_key[1119]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1119]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1119]               =   1'b0;
assign   tb_i_rf_static_encrypt[1119]          =   1'b1;
assign   tb_i_clear_fault_flags[1119]          =   1'b0;
assign   tb_i_rf_static_aad_length[1119]       =   64'h0000000000000100;
assign   tb_i_aad[1119]                        =   tb_i_aad[1118];
assign   tb_i_rf_static_plaintext_length[1119] =   64'h0000000000000280;
assign   tb_i_plaintext[1119]                  =   tb_i_plaintext[1118];
assign   tb_o_valid[1119]                      =   1'b0;
assign   tb_o_sop[1119]                        =   1'b0;
assign   tb_o_ciphertext[1119]                 =   tb_o_ciphertext[1118];
assign   tb_o_tag_ready[1119]                  =   1'b1;
assign   tb_o_tag[1119]                        =   128'hb4a1b3d8763ca30d7bbd2894b60718c6;

// CLK no. 1120/1240
// *************************************************
assign   tb_i_valid[1120]                      =   1'b0;
assign   tb_i_reset[1120]                      =   1'b0;
assign   tb_i_sop[1120]                        =   1'b0;
assign   tb_i_key_update[1120]                 =   1'b0;
assign   tb_i_key[1120]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1120]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1120]               =   1'b0;
assign   tb_i_rf_static_encrypt[1120]          =   1'b1;
assign   tb_i_clear_fault_flags[1120]          =   1'b0;
assign   tb_i_rf_static_aad_length[1120]       =   64'h0000000000000100;
assign   tb_i_aad[1120]                        =   tb_i_aad[1119];
assign   tb_i_rf_static_plaintext_length[1120] =   64'h0000000000000280;
assign   tb_i_plaintext[1120]                  =   tb_i_plaintext[1119];
assign   tb_o_valid[1120]                      =   1'b0;
assign   tb_o_sop[1120]                        =   1'b0;
assign   tb_o_ciphertext[1120]                 =   tb_o_ciphertext[1119];
assign   tb_o_tag_ready[1120]                  =   1'b0;
assign   tb_o_tag[1120]                        =   tb_o_tag[1119];

// CLK no. 1121/1240
// *************************************************
assign   tb_i_valid[1121]                      =   1'b0;
assign   tb_i_reset[1121]                      =   1'b0;
assign   tb_i_sop[1121]                        =   1'b0;
assign   tb_i_key_update[1121]                 =   1'b0;
assign   tb_i_key[1121]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1121]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1121]               =   1'b0;
assign   tb_i_rf_static_encrypt[1121]          =   1'b1;
assign   tb_i_clear_fault_flags[1121]          =   1'b0;
assign   tb_i_rf_static_aad_length[1121]       =   64'h0000000000000100;
assign   tb_i_aad[1121]                        =   tb_i_aad[1120];
assign   tb_i_rf_static_plaintext_length[1121] =   64'h0000000000000280;
assign   tb_i_plaintext[1121]                  =   tb_i_plaintext[1120];
assign   tb_o_valid[1121]                      =   1'b0;
assign   tb_o_sop[1121]                        =   1'b0;
assign   tb_o_ciphertext[1121]                 =   tb_o_ciphertext[1120];
assign   tb_o_tag_ready[1121]                  =   1'b0;
assign   tb_o_tag[1121]                        =   tb_o_tag[1120];

// CLK no. 1122/1240
// *************************************************
assign   tb_i_valid[1122]                      =   1'b0;
assign   tb_i_reset[1122]                      =   1'b0;
assign   tb_i_sop[1122]                        =   1'b1;
assign   tb_i_key_update[1122]                 =   1'b0;
assign   tb_i_key[1122]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1122]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1122]               =   1'b0;
assign   tb_i_rf_static_encrypt[1122]          =   1'b1;
assign   tb_i_clear_fault_flags[1122]          =   1'b0;
assign   tb_i_rf_static_aad_length[1122]       =   64'h0000000000000100;
assign   tb_i_aad[1122]                        =   tb_i_aad[1121];
assign   tb_i_rf_static_plaintext_length[1122] =   64'h0000000000000280;
assign   tb_i_plaintext[1122]                  =   tb_i_plaintext[1121];
assign   tb_o_valid[1122]                      =   1'b0;
assign   tb_o_sop[1122]                        =   1'b0;
assign   tb_o_ciphertext[1122]                 =   tb_o_ciphertext[1121];
assign   tb_o_tag_ready[1122]                  =   1'b0;
assign   tb_o_tag[1122]                        =   tb_o_tag[1121];

// CLK no. 1123/1240
// *************************************************
assign   tb_i_valid[1123]                      =   1'b1;
assign   tb_i_reset[1123]                      =   1'b0;
assign   tb_i_sop[1123]                        =   1'b0;
assign   tb_i_key_update[1123]                 =   1'b0;
assign   tb_i_key[1123]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1123]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1123]               =   1'b0;
assign   tb_i_rf_static_encrypt[1123]          =   1'b1;
assign   tb_i_clear_fault_flags[1123]          =   1'b0;
assign   tb_i_rf_static_aad_length[1123]       =   64'h0000000000000100;
assign   tb_i_aad[1123]                        =   256'h990ee47fb832543e894038d5b2a76619a9b399699824d6861a04c6608c039d06;
assign   tb_i_rf_static_plaintext_length[1123] =   64'h0000000000000280;
assign   tb_i_plaintext[1123]                  =   tb_i_plaintext[1122];
assign   tb_o_valid[1123]                      =   1'b0;
assign   tb_o_sop[1123]                        =   1'b0;
assign   tb_o_ciphertext[1123]                 =   tb_o_ciphertext[1122];
assign   tb_o_tag_ready[1123]                  =   1'b0;
assign   tb_o_tag[1123]                        =   tb_o_tag[1122];

// CLK no. 1124/1240
// *************************************************
assign   tb_i_valid[1124]                      =   1'b1;
assign   tb_i_reset[1124]                      =   1'b0;
assign   tb_i_sop[1124]                        =   1'b0;
assign   tb_i_key_update[1124]                 =   1'b0;
assign   tb_i_key[1124]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1124]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1124]               =   1'b0;
assign   tb_i_rf_static_encrypt[1124]          =   1'b1;
assign   tb_i_clear_fault_flags[1124]          =   1'b0;
assign   tb_i_rf_static_aad_length[1124]       =   64'h0000000000000100;
assign   tb_i_aad[1124]                        =   tb_i_aad[1123];
assign   tb_i_rf_static_plaintext_length[1124] =   64'h0000000000000280;
assign   tb_i_plaintext[1124]                  =   256'ha4b1f15b1c2d1ef4b8f18635f25b0af3a55354ff812d51d34f8fad0cc936b048;
assign   tb_o_valid[1124]                      =   1'b0;
assign   tb_o_sop[1124]                        =   1'b0;
assign   tb_o_ciphertext[1124]                 =   tb_o_ciphertext[1123];
assign   tb_o_tag_ready[1124]                  =   1'b0;
assign   tb_o_tag[1124]                        =   tb_o_tag[1123];

// CLK no. 1125/1240
// *************************************************
assign   tb_i_valid[1125]                      =   1'b1;
assign   tb_i_reset[1125]                      =   1'b0;
assign   tb_i_sop[1125]                        =   1'b0;
assign   tb_i_key_update[1125]                 =   1'b0;
assign   tb_i_key[1125]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1125]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1125]               =   1'b0;
assign   tb_i_rf_static_encrypt[1125]          =   1'b1;
assign   tb_i_clear_fault_flags[1125]          =   1'b0;
assign   tb_i_rf_static_aad_length[1125]       =   64'h0000000000000100;
assign   tb_i_aad[1125]                        =   tb_i_aad[1124];
assign   tb_i_rf_static_plaintext_length[1125] =   64'h0000000000000280;
assign   tb_i_plaintext[1125]                  =   256'h7059bd045aaff8ff4ef882e79873ac58a061ccff534307664edf592502a2b828;
assign   tb_o_valid[1125]                      =   1'b0;
assign   tb_o_sop[1125]                        =   1'b0;
assign   tb_o_ciphertext[1125]                 =   tb_o_ciphertext[1124];
assign   tb_o_tag_ready[1125]                  =   1'b0;
assign   tb_o_tag[1125]                        =   tb_o_tag[1124];

// CLK no. 1126/1240
// *************************************************
assign   tb_i_valid[1126]                      =   1'b1;
assign   tb_i_reset[1126]                      =   1'b0;
assign   tb_i_sop[1126]                        =   1'b0;
assign   tb_i_key_update[1126]                 =   1'b0;
assign   tb_i_key[1126]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1126]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1126]               =   1'b0;
assign   tb_i_rf_static_encrypt[1126]          =   1'b1;
assign   tb_i_clear_fault_flags[1126]          =   1'b0;
assign   tb_i_rf_static_aad_length[1126]       =   64'h0000000000000100;
assign   tb_i_aad[1126]                        =   tb_i_aad[1125];
assign   tb_i_rf_static_plaintext_length[1126] =   64'h0000000000000280;
assign   tb_i_plaintext[1126]                  =   256'hf6932830ae7fc0ac41a5b5bcf5c87d08;
assign   tb_o_valid[1126]                      =   1'b0;
assign   tb_o_sop[1126]                        =   1'b0;
assign   tb_o_ciphertext[1126]                 =   tb_o_ciphertext[1125];
assign   tb_o_tag_ready[1126]                  =   1'b0;
assign   tb_o_tag[1126]                        =   tb_o_tag[1125];

// CLK no. 1127/1240
// *************************************************
assign   tb_i_valid[1127]                      =   1'b0;
assign   tb_i_reset[1127]                      =   1'b0;
assign   tb_i_sop[1127]                        =   1'b0;
assign   tb_i_key_update[1127]                 =   1'b0;
assign   tb_i_key[1127]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1127]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1127]               =   1'b0;
assign   tb_i_rf_static_encrypt[1127]          =   1'b1;
assign   tb_i_clear_fault_flags[1127]          =   1'b0;
assign   tb_i_rf_static_aad_length[1127]       =   64'h0000000000000100;
assign   tb_i_aad[1127]                        =   tb_i_aad[1126];
assign   tb_i_rf_static_plaintext_length[1127] =   64'h0000000000000280;
assign   tb_i_plaintext[1127]                  =   tb_i_plaintext[1126];
assign   tb_o_valid[1127]                      =   1'b0;
assign   tb_o_sop[1127]                        =   1'b0;
assign   tb_o_ciphertext[1127]                 =   tb_o_ciphertext[1126];
assign   tb_o_tag_ready[1127]                  =   1'b0;
assign   tb_o_tag[1127]                        =   tb_o_tag[1126];

// CLK no. 1128/1240
// *************************************************
assign   tb_i_valid[1128]                      =   1'b0;
assign   tb_i_reset[1128]                      =   1'b0;
assign   tb_i_sop[1128]                        =   1'b0;
assign   tb_i_key_update[1128]                 =   1'b0;
assign   tb_i_key[1128]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1128]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1128]               =   1'b0;
assign   tb_i_rf_static_encrypt[1128]          =   1'b1;
assign   tb_i_clear_fault_flags[1128]          =   1'b0;
assign   tb_i_rf_static_aad_length[1128]       =   64'h0000000000000100;
assign   tb_i_aad[1128]                        =   tb_i_aad[1127];
assign   tb_i_rf_static_plaintext_length[1128] =   64'h0000000000000280;
assign   tb_i_plaintext[1128]                  =   tb_i_plaintext[1127];
assign   tb_o_valid[1128]                      =   1'b0;
assign   tb_o_sop[1128]                        =   1'b0;
assign   tb_o_ciphertext[1128]                 =   tb_o_ciphertext[1127];
assign   tb_o_tag_ready[1128]                  =   1'b0;
assign   tb_o_tag[1128]                        =   tb_o_tag[1127];

// CLK no. 1129/1240
// *************************************************
assign   tb_i_valid[1129]                      =   1'b0;
assign   tb_i_reset[1129]                      =   1'b0;
assign   tb_i_sop[1129]                        =   1'b0;
assign   tb_i_key_update[1129]                 =   1'b0;
assign   tb_i_key[1129]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1129]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1129]               =   1'b0;
assign   tb_i_rf_static_encrypt[1129]          =   1'b1;
assign   tb_i_clear_fault_flags[1129]          =   1'b0;
assign   tb_i_rf_static_aad_length[1129]       =   64'h0000000000000100;
assign   tb_i_aad[1129]                        =   tb_i_aad[1128];
assign   tb_i_rf_static_plaintext_length[1129] =   64'h0000000000000280;
assign   tb_i_plaintext[1129]                  =   tb_i_plaintext[1128];
assign   tb_o_valid[1129]                      =   1'b0;
assign   tb_o_sop[1129]                        =   1'b0;
assign   tb_o_ciphertext[1129]                 =   tb_o_ciphertext[1128];
assign   tb_o_tag_ready[1129]                  =   1'b0;
assign   tb_o_tag[1129]                        =   tb_o_tag[1128];

// CLK no. 1130/1240
// *************************************************
assign   tb_i_valid[1130]                      =   1'b0;
assign   tb_i_reset[1130]                      =   1'b0;
assign   tb_i_sop[1130]                        =   1'b0;
assign   tb_i_key_update[1130]                 =   1'b0;
assign   tb_i_key[1130]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1130]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1130]               =   1'b0;
assign   tb_i_rf_static_encrypt[1130]          =   1'b1;
assign   tb_i_clear_fault_flags[1130]          =   1'b0;
assign   tb_i_rf_static_aad_length[1130]       =   64'h0000000000000100;
assign   tb_i_aad[1130]                        =   tb_i_aad[1129];
assign   tb_i_rf_static_plaintext_length[1130] =   64'h0000000000000280;
assign   tb_i_plaintext[1130]                  =   tb_i_plaintext[1129];
assign   tb_o_valid[1130]                      =   1'b0;
assign   tb_o_sop[1130]                        =   1'b0;
assign   tb_o_ciphertext[1130]                 =   tb_o_ciphertext[1129];
assign   tb_o_tag_ready[1130]                  =   1'b0;
assign   tb_o_tag[1130]                        =   tb_o_tag[1129];

// CLK no. 1131/1240
// *************************************************
assign   tb_i_valid[1131]                      =   1'b0;
assign   tb_i_reset[1131]                      =   1'b0;
assign   tb_i_sop[1131]                        =   1'b0;
assign   tb_i_key_update[1131]                 =   1'b0;
assign   tb_i_key[1131]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1131]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1131]               =   1'b0;
assign   tb_i_rf_static_encrypt[1131]          =   1'b1;
assign   tb_i_clear_fault_flags[1131]          =   1'b0;
assign   tb_i_rf_static_aad_length[1131]       =   64'h0000000000000100;
assign   tb_i_aad[1131]                        =   tb_i_aad[1130];
assign   tb_i_rf_static_plaintext_length[1131] =   64'h0000000000000280;
assign   tb_i_plaintext[1131]                  =   tb_i_plaintext[1130];
assign   tb_o_valid[1131]                      =   1'b0;
assign   tb_o_sop[1131]                        =   1'b0;
assign   tb_o_ciphertext[1131]                 =   tb_o_ciphertext[1130];
assign   tb_o_tag_ready[1131]                  =   1'b0;
assign   tb_o_tag[1131]                        =   tb_o_tag[1130];

// CLK no. 1132/1240
// *************************************************
assign   tb_i_valid[1132]                      =   1'b0;
assign   tb_i_reset[1132]                      =   1'b0;
assign   tb_i_sop[1132]                        =   1'b0;
assign   tb_i_key_update[1132]                 =   1'b0;
assign   tb_i_key[1132]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1132]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1132]               =   1'b0;
assign   tb_i_rf_static_encrypt[1132]          =   1'b1;
assign   tb_i_clear_fault_flags[1132]          =   1'b0;
assign   tb_i_rf_static_aad_length[1132]       =   64'h0000000000000100;
assign   tb_i_aad[1132]                        =   tb_i_aad[1131];
assign   tb_i_rf_static_plaintext_length[1132] =   64'h0000000000000280;
assign   tb_i_plaintext[1132]                  =   tb_i_plaintext[1131];
assign   tb_o_valid[1132]                      =   1'b0;
assign   tb_o_sop[1132]                        =   1'b0;
assign   tb_o_ciphertext[1132]                 =   tb_o_ciphertext[1131];
assign   tb_o_tag_ready[1132]                  =   1'b0;
assign   tb_o_tag[1132]                        =   tb_o_tag[1131];

// CLK no. 1133/1240
// *************************************************
assign   tb_i_valid[1133]                      =   1'b0;
assign   tb_i_reset[1133]                      =   1'b0;
assign   tb_i_sop[1133]                        =   1'b0;
assign   tb_i_key_update[1133]                 =   1'b0;
assign   tb_i_key[1133]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1133]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1133]               =   1'b0;
assign   tb_i_rf_static_encrypt[1133]          =   1'b1;
assign   tb_i_clear_fault_flags[1133]          =   1'b0;
assign   tb_i_rf_static_aad_length[1133]       =   64'h0000000000000100;
assign   tb_i_aad[1133]                        =   tb_i_aad[1132];
assign   tb_i_rf_static_plaintext_length[1133] =   64'h0000000000000280;
assign   tb_i_plaintext[1133]                  =   tb_i_plaintext[1132];
assign   tb_o_valid[1133]                      =   1'b0;
assign   tb_o_sop[1133]                        =   1'b0;
assign   tb_o_ciphertext[1133]                 =   tb_o_ciphertext[1132];
assign   tb_o_tag_ready[1133]                  =   1'b0;
assign   tb_o_tag[1133]                        =   tb_o_tag[1132];

// CLK no. 1134/1240
// *************************************************
assign   tb_i_valid[1134]                      =   1'b0;
assign   tb_i_reset[1134]                      =   1'b0;
assign   tb_i_sop[1134]                        =   1'b0;
assign   tb_i_key_update[1134]                 =   1'b0;
assign   tb_i_key[1134]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1134]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1134]               =   1'b0;
assign   tb_i_rf_static_encrypt[1134]          =   1'b1;
assign   tb_i_clear_fault_flags[1134]          =   1'b0;
assign   tb_i_rf_static_aad_length[1134]       =   64'h0000000000000100;
assign   tb_i_aad[1134]                        =   tb_i_aad[1133];
assign   tb_i_rf_static_plaintext_length[1134] =   64'h0000000000000280;
assign   tb_i_plaintext[1134]                  =   tb_i_plaintext[1133];
assign   tb_o_valid[1134]                      =   1'b0;
assign   tb_o_sop[1134]                        =   1'b0;
assign   tb_o_ciphertext[1134]                 =   tb_o_ciphertext[1133];
assign   tb_o_tag_ready[1134]                  =   1'b0;
assign   tb_o_tag[1134]                        =   tb_o_tag[1133];

// CLK no. 1135/1240
// *************************************************
assign   tb_i_valid[1135]                      =   1'b0;
assign   tb_i_reset[1135]                      =   1'b0;
assign   tb_i_sop[1135]                        =   1'b0;
assign   tb_i_key_update[1135]                 =   1'b0;
assign   tb_i_key[1135]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1135]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1135]               =   1'b0;
assign   tb_i_rf_static_encrypt[1135]          =   1'b1;
assign   tb_i_clear_fault_flags[1135]          =   1'b0;
assign   tb_i_rf_static_aad_length[1135]       =   64'h0000000000000100;
assign   tb_i_aad[1135]                        =   tb_i_aad[1134];
assign   tb_i_rf_static_plaintext_length[1135] =   64'h0000000000000280;
assign   tb_i_plaintext[1135]                  =   tb_i_plaintext[1134];
assign   tb_o_valid[1135]                      =   1'b0;
assign   tb_o_sop[1135]                        =   1'b0;
assign   tb_o_ciphertext[1135]                 =   tb_o_ciphertext[1134];
assign   tb_o_tag_ready[1135]                  =   1'b0;
assign   tb_o_tag[1135]                        =   tb_o_tag[1134];

// CLK no. 1136/1240
// *************************************************
assign   tb_i_valid[1136]                      =   1'b0;
assign   tb_i_reset[1136]                      =   1'b0;
assign   tb_i_sop[1136]                        =   1'b0;
assign   tb_i_key_update[1136]                 =   1'b0;
assign   tb_i_key[1136]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1136]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1136]               =   1'b0;
assign   tb_i_rf_static_encrypt[1136]          =   1'b1;
assign   tb_i_clear_fault_flags[1136]          =   1'b0;
assign   tb_i_rf_static_aad_length[1136]       =   64'h0000000000000100;
assign   tb_i_aad[1136]                        =   tb_i_aad[1135];
assign   tb_i_rf_static_plaintext_length[1136] =   64'h0000000000000280;
assign   tb_i_plaintext[1136]                  =   tb_i_plaintext[1135];
assign   tb_o_valid[1136]                      =   1'b0;
assign   tb_o_sop[1136]                        =   1'b0;
assign   tb_o_ciphertext[1136]                 =   tb_o_ciphertext[1135];
assign   tb_o_tag_ready[1136]                  =   1'b0;
assign   tb_o_tag[1136]                        =   tb_o_tag[1135];

// CLK no. 1137/1240
// *************************************************
assign   tb_i_valid[1137]                      =   1'b0;
assign   tb_i_reset[1137]                      =   1'b0;
assign   tb_i_sop[1137]                        =   1'b0;
assign   tb_i_key_update[1137]                 =   1'b0;
assign   tb_i_key[1137]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1137]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1137]               =   1'b0;
assign   tb_i_rf_static_encrypt[1137]          =   1'b1;
assign   tb_i_clear_fault_flags[1137]          =   1'b0;
assign   tb_i_rf_static_aad_length[1137]       =   64'h0000000000000100;
assign   tb_i_aad[1137]                        =   tb_i_aad[1136];
assign   tb_i_rf_static_plaintext_length[1137] =   64'h0000000000000280;
assign   tb_i_plaintext[1137]                  =   tb_i_plaintext[1136];
assign   tb_o_valid[1137]                      =   1'b0;
assign   tb_o_sop[1137]                        =   1'b0;
assign   tb_o_ciphertext[1137]                 =   tb_o_ciphertext[1136];
assign   tb_o_tag_ready[1137]                  =   1'b0;
assign   tb_o_tag[1137]                        =   tb_o_tag[1136];

// CLK no. 1138/1240
// *************************************************
assign   tb_i_valid[1138]                      =   1'b0;
assign   tb_i_reset[1138]                      =   1'b0;
assign   tb_i_sop[1138]                        =   1'b0;
assign   tb_i_key_update[1138]                 =   1'b0;
assign   tb_i_key[1138]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1138]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1138]               =   1'b0;
assign   tb_i_rf_static_encrypt[1138]          =   1'b1;
assign   tb_i_clear_fault_flags[1138]          =   1'b0;
assign   tb_i_rf_static_aad_length[1138]       =   64'h0000000000000100;
assign   tb_i_aad[1138]                        =   tb_i_aad[1137];
assign   tb_i_rf_static_plaintext_length[1138] =   64'h0000000000000280;
assign   tb_i_plaintext[1138]                  =   tb_i_plaintext[1137];
assign   tb_o_valid[1138]                      =   1'b0;
assign   tb_o_sop[1138]                        =   1'b0;
assign   tb_o_ciphertext[1138]                 =   tb_o_ciphertext[1137];
assign   tb_o_tag_ready[1138]                  =   1'b0;
assign   tb_o_tag[1138]                        =   tb_o_tag[1137];

// CLK no. 1139/1240
// *************************************************
assign   tb_i_valid[1139]                      =   1'b0;
assign   tb_i_reset[1139]                      =   1'b0;
assign   tb_i_sop[1139]                        =   1'b0;
assign   tb_i_key_update[1139]                 =   1'b0;
assign   tb_i_key[1139]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1139]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1139]               =   1'b0;
assign   tb_i_rf_static_encrypt[1139]          =   1'b1;
assign   tb_i_clear_fault_flags[1139]          =   1'b0;
assign   tb_i_rf_static_aad_length[1139]       =   64'h0000000000000100;
assign   tb_i_aad[1139]                        =   tb_i_aad[1138];
assign   tb_i_rf_static_plaintext_length[1139] =   64'h0000000000000280;
assign   tb_i_plaintext[1139]                  =   tb_i_plaintext[1138];
assign   tb_o_valid[1139]                      =   1'b0;
assign   tb_o_sop[1139]                        =   1'b0;
assign   tb_o_ciphertext[1139]                 =   tb_o_ciphertext[1138];
assign   tb_o_tag_ready[1139]                  =   1'b0;
assign   tb_o_tag[1139]                        =   tb_o_tag[1138];

// CLK no. 1140/1240
// *************************************************
assign   tb_i_valid[1140]                      =   1'b0;
assign   tb_i_reset[1140]                      =   1'b0;
assign   tb_i_sop[1140]                        =   1'b0;
assign   tb_i_key_update[1140]                 =   1'b0;
assign   tb_i_key[1140]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1140]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1140]               =   1'b0;
assign   tb_i_rf_static_encrypt[1140]          =   1'b1;
assign   tb_i_clear_fault_flags[1140]          =   1'b0;
assign   tb_i_rf_static_aad_length[1140]       =   64'h0000000000000100;
assign   tb_i_aad[1140]                        =   tb_i_aad[1139];
assign   tb_i_rf_static_plaintext_length[1140] =   64'h0000000000000280;
assign   tb_i_plaintext[1140]                  =   tb_i_plaintext[1139];
assign   tb_o_valid[1140]                      =   1'b0;
assign   tb_o_sop[1140]                        =   1'b0;
assign   tb_o_ciphertext[1140]                 =   tb_o_ciphertext[1139];
assign   tb_o_tag_ready[1140]                  =   1'b0;
assign   tb_o_tag[1140]                        =   tb_o_tag[1139];

// CLK no. 1141/1240
// *************************************************
assign   tb_i_valid[1141]                      =   1'b0;
assign   tb_i_reset[1141]                      =   1'b0;
assign   tb_i_sop[1141]                        =   1'b0;
assign   tb_i_key_update[1141]                 =   1'b0;
assign   tb_i_key[1141]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1141]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1141]               =   1'b0;
assign   tb_i_rf_static_encrypt[1141]          =   1'b1;
assign   tb_i_clear_fault_flags[1141]          =   1'b0;
assign   tb_i_rf_static_aad_length[1141]       =   64'h0000000000000100;
assign   tb_i_aad[1141]                        =   tb_i_aad[1140];
assign   tb_i_rf_static_plaintext_length[1141] =   64'h0000000000000280;
assign   tb_i_plaintext[1141]                  =   tb_i_plaintext[1140];
assign   tb_o_valid[1141]                      =   1'b0;
assign   tb_o_sop[1141]                        =   1'b0;
assign   tb_o_ciphertext[1141]                 =   tb_o_ciphertext[1140];
assign   tb_o_tag_ready[1141]                  =   1'b0;
assign   tb_o_tag[1141]                        =   tb_o_tag[1140];

// CLK no. 1142/1240
// *************************************************
assign   tb_i_valid[1142]                      =   1'b0;
assign   tb_i_reset[1142]                      =   1'b0;
assign   tb_i_sop[1142]                        =   1'b0;
assign   tb_i_key_update[1142]                 =   1'b0;
assign   tb_i_key[1142]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1142]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1142]               =   1'b0;
assign   tb_i_rf_static_encrypt[1142]          =   1'b1;
assign   tb_i_clear_fault_flags[1142]          =   1'b0;
assign   tb_i_rf_static_aad_length[1142]       =   64'h0000000000000100;
assign   tb_i_aad[1142]                        =   tb_i_aad[1141];
assign   tb_i_rf_static_plaintext_length[1142] =   64'h0000000000000280;
assign   tb_i_plaintext[1142]                  =   tb_i_plaintext[1141];
assign   tb_o_valid[1142]                      =   1'b0;
assign   tb_o_sop[1142]                        =   1'b0;
assign   tb_o_ciphertext[1142]                 =   tb_o_ciphertext[1141];
assign   tb_o_tag_ready[1142]                  =   1'b0;
assign   tb_o_tag[1142]                        =   tb_o_tag[1141];

// CLK no. 1143/1240
// *************************************************
assign   tb_i_valid[1143]                      =   1'b0;
assign   tb_i_reset[1143]                      =   1'b0;
assign   tb_i_sop[1143]                        =   1'b0;
assign   tb_i_key_update[1143]                 =   1'b0;
assign   tb_i_key[1143]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1143]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1143]               =   1'b0;
assign   tb_i_rf_static_encrypt[1143]          =   1'b1;
assign   tb_i_clear_fault_flags[1143]          =   1'b0;
assign   tb_i_rf_static_aad_length[1143]       =   64'h0000000000000100;
assign   tb_i_aad[1143]                        =   tb_i_aad[1142];
assign   tb_i_rf_static_plaintext_length[1143] =   64'h0000000000000280;
assign   tb_i_plaintext[1143]                  =   tb_i_plaintext[1142];
assign   tb_o_valid[1143]                      =   1'b0;
assign   tb_o_sop[1143]                        =   1'b0;
assign   tb_o_ciphertext[1143]                 =   tb_o_ciphertext[1142];
assign   tb_o_tag_ready[1143]                  =   1'b0;
assign   tb_o_tag[1143]                        =   tb_o_tag[1142];

// CLK no. 1144/1240
// *************************************************
assign   tb_i_valid[1144]                      =   1'b0;
assign   tb_i_reset[1144]                      =   1'b0;
assign   tb_i_sop[1144]                        =   1'b0;
assign   tb_i_key_update[1144]                 =   1'b0;
assign   tb_i_key[1144]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1144]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1144]               =   1'b0;
assign   tb_i_rf_static_encrypt[1144]          =   1'b1;
assign   tb_i_clear_fault_flags[1144]          =   1'b0;
assign   tb_i_rf_static_aad_length[1144]       =   64'h0000000000000100;
assign   tb_i_aad[1144]                        =   tb_i_aad[1143];
assign   tb_i_rf_static_plaintext_length[1144] =   64'h0000000000000280;
assign   tb_i_plaintext[1144]                  =   tb_i_plaintext[1143];
assign   tb_o_valid[1144]                      =   1'b0;
assign   tb_o_sop[1144]                        =   1'b0;
assign   tb_o_ciphertext[1144]                 =   tb_o_ciphertext[1143];
assign   tb_o_tag_ready[1144]                  =   1'b0;
assign   tb_o_tag[1144]                        =   tb_o_tag[1143];

// CLK no. 1145/1240
// *************************************************
assign   tb_i_valid[1145]                      =   1'b0;
assign   tb_i_reset[1145]                      =   1'b0;
assign   tb_i_sop[1145]                        =   1'b0;
assign   tb_i_key_update[1145]                 =   1'b0;
assign   tb_i_key[1145]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1145]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1145]               =   1'b0;
assign   tb_i_rf_static_encrypt[1145]          =   1'b1;
assign   tb_i_clear_fault_flags[1145]          =   1'b0;
assign   tb_i_rf_static_aad_length[1145]       =   64'h0000000000000100;
assign   tb_i_aad[1145]                        =   tb_i_aad[1144];
assign   tb_i_rf_static_plaintext_length[1145] =   64'h0000000000000280;
assign   tb_i_plaintext[1145]                  =   tb_i_plaintext[1144];
assign   tb_o_valid[1145]                      =   1'b0;
assign   tb_o_sop[1145]                        =   1'b0;
assign   tb_o_ciphertext[1145]                 =   tb_o_ciphertext[1144];
assign   tb_o_tag_ready[1145]                  =   1'b0;
assign   tb_o_tag[1145]                        =   tb_o_tag[1144];

// CLK no. 1146/1240
// *************************************************
assign   tb_i_valid[1146]                      =   1'b0;
assign   tb_i_reset[1146]                      =   1'b0;
assign   tb_i_sop[1146]                        =   1'b0;
assign   tb_i_key_update[1146]                 =   1'b0;
assign   tb_i_key[1146]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1146]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1146]               =   1'b0;
assign   tb_i_rf_static_encrypt[1146]          =   1'b1;
assign   tb_i_clear_fault_flags[1146]          =   1'b0;
assign   tb_i_rf_static_aad_length[1146]       =   64'h0000000000000100;
assign   tb_i_aad[1146]                        =   tb_i_aad[1145];
assign   tb_i_rf_static_plaintext_length[1146] =   64'h0000000000000280;
assign   tb_i_plaintext[1146]                  =   tb_i_plaintext[1145];
assign   tb_o_valid[1146]                      =   1'b0;
assign   tb_o_sop[1146]                        =   1'b0;
assign   tb_o_ciphertext[1146]                 =   tb_o_ciphertext[1145];
assign   tb_o_tag_ready[1146]                  =   1'b0;
assign   tb_o_tag[1146]                        =   tb_o_tag[1145];

// CLK no. 1147/1240
// *************************************************
assign   tb_i_valid[1147]                      =   1'b0;
assign   tb_i_reset[1147]                      =   1'b0;
assign   tb_i_sop[1147]                        =   1'b0;
assign   tb_i_key_update[1147]                 =   1'b0;
assign   tb_i_key[1147]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1147]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1147]               =   1'b0;
assign   tb_i_rf_static_encrypt[1147]          =   1'b1;
assign   tb_i_clear_fault_flags[1147]          =   1'b0;
assign   tb_i_rf_static_aad_length[1147]       =   64'h0000000000000100;
assign   tb_i_aad[1147]                        =   tb_i_aad[1146];
assign   tb_i_rf_static_plaintext_length[1147] =   64'h0000000000000280;
assign   tb_i_plaintext[1147]                  =   tb_i_plaintext[1146];
assign   tb_o_valid[1147]                      =   1'b0;
assign   tb_o_sop[1147]                        =   1'b0;
assign   tb_o_ciphertext[1147]                 =   tb_o_ciphertext[1146];
assign   tb_o_tag_ready[1147]                  =   1'b0;
assign   tb_o_tag[1147]                        =   tb_o_tag[1146];

// CLK no. 1148/1240
// *************************************************
assign   tb_i_valid[1148]                      =   1'b0;
assign   tb_i_reset[1148]                      =   1'b0;
assign   tb_i_sop[1148]                        =   1'b0;
assign   tb_i_key_update[1148]                 =   1'b0;
assign   tb_i_key[1148]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1148]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1148]               =   1'b0;
assign   tb_i_rf_static_encrypt[1148]          =   1'b1;
assign   tb_i_clear_fault_flags[1148]          =   1'b0;
assign   tb_i_rf_static_aad_length[1148]       =   64'h0000000000000100;
assign   tb_i_aad[1148]                        =   tb_i_aad[1147];
assign   tb_i_rf_static_plaintext_length[1148] =   64'h0000000000000280;
assign   tb_i_plaintext[1148]                  =   tb_i_plaintext[1147];
assign   tb_o_valid[1148]                      =   1'b0;
assign   tb_o_sop[1148]                        =   1'b0;
assign   tb_o_ciphertext[1148]                 =   tb_o_ciphertext[1147];
assign   tb_o_tag_ready[1148]                  =   1'b0;
assign   tb_o_tag[1148]                        =   tb_o_tag[1147];

// CLK no. 1149/1240
// *************************************************
assign   tb_i_valid[1149]                      =   1'b0;
assign   tb_i_reset[1149]                      =   1'b0;
assign   tb_i_sop[1149]                        =   1'b0;
assign   tb_i_key_update[1149]                 =   1'b0;
assign   tb_i_key[1149]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1149]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1149]               =   1'b0;
assign   tb_i_rf_static_encrypt[1149]          =   1'b1;
assign   tb_i_clear_fault_flags[1149]          =   1'b0;
assign   tb_i_rf_static_aad_length[1149]       =   64'h0000000000000100;
assign   tb_i_aad[1149]                        =   tb_i_aad[1148];
assign   tb_i_rf_static_plaintext_length[1149] =   64'h0000000000000280;
assign   tb_i_plaintext[1149]                  =   tb_i_plaintext[1148];
assign   tb_o_valid[1149]                      =   1'b0;
assign   tb_o_sop[1149]                        =   1'b0;
assign   tb_o_ciphertext[1149]                 =   tb_o_ciphertext[1148];
assign   tb_o_tag_ready[1149]                  =   1'b0;
assign   tb_o_tag[1149]                        =   tb_o_tag[1148];

// CLK no. 1150/1240
// *************************************************
assign   tb_i_valid[1150]                      =   1'b0;
assign   tb_i_reset[1150]                      =   1'b0;
assign   tb_i_sop[1150]                        =   1'b0;
assign   tb_i_key_update[1150]                 =   1'b0;
assign   tb_i_key[1150]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1150]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1150]               =   1'b0;
assign   tb_i_rf_static_encrypt[1150]          =   1'b1;
assign   tb_i_clear_fault_flags[1150]          =   1'b0;
assign   tb_i_rf_static_aad_length[1150]       =   64'h0000000000000100;
assign   tb_i_aad[1150]                        =   tb_i_aad[1149];
assign   tb_i_rf_static_plaintext_length[1150] =   64'h0000000000000280;
assign   tb_i_plaintext[1150]                  =   tb_i_plaintext[1149];
assign   tb_o_valid[1150]                      =   1'b0;
assign   tb_o_sop[1150]                        =   1'b0;
assign   tb_o_ciphertext[1150]                 =   tb_o_ciphertext[1149];
assign   tb_o_tag_ready[1150]                  =   1'b0;
assign   tb_o_tag[1150]                        =   tb_o_tag[1149];

// CLK no. 1151/1240
// *************************************************
assign   tb_i_valid[1151]                      =   1'b0;
assign   tb_i_reset[1151]                      =   1'b0;
assign   tb_i_sop[1151]                        =   1'b0;
assign   tb_i_key_update[1151]                 =   1'b0;
assign   tb_i_key[1151]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1151]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1151]               =   1'b0;
assign   tb_i_rf_static_encrypt[1151]          =   1'b1;
assign   tb_i_clear_fault_flags[1151]          =   1'b0;
assign   tb_i_rf_static_aad_length[1151]       =   64'h0000000000000100;
assign   tb_i_aad[1151]                        =   tb_i_aad[1150];
assign   tb_i_rf_static_plaintext_length[1151] =   64'h0000000000000280;
assign   tb_i_plaintext[1151]                  =   tb_i_plaintext[1150];
assign   tb_o_valid[1151]                      =   1'b0;
assign   tb_o_sop[1151]                        =   1'b0;
assign   tb_o_ciphertext[1151]                 =   tb_o_ciphertext[1150];
assign   tb_o_tag_ready[1151]                  =   1'b0;
assign   tb_o_tag[1151]                        =   tb_o_tag[1150];

// CLK no. 1152/1240
// *************************************************
assign   tb_i_valid[1152]                      =   1'b0;
assign   tb_i_reset[1152]                      =   1'b0;
assign   tb_i_sop[1152]                        =   1'b0;
assign   tb_i_key_update[1152]                 =   1'b0;
assign   tb_i_key[1152]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1152]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1152]               =   1'b0;
assign   tb_i_rf_static_encrypt[1152]          =   1'b1;
assign   tb_i_clear_fault_flags[1152]          =   1'b0;
assign   tb_i_rf_static_aad_length[1152]       =   64'h0000000000000100;
assign   tb_i_aad[1152]                        =   tb_i_aad[1151];
assign   tb_i_rf_static_plaintext_length[1152] =   64'h0000000000000280;
assign   tb_i_plaintext[1152]                  =   tb_i_plaintext[1151];
assign   tb_o_valid[1152]                      =   1'b0;
assign   tb_o_sop[1152]                        =   1'b0;
assign   tb_o_ciphertext[1152]                 =   tb_o_ciphertext[1151];
assign   tb_o_tag_ready[1152]                  =   1'b0;
assign   tb_o_tag[1152]                        =   tb_o_tag[1151];

// CLK no. 1153/1240
// *************************************************
assign   tb_i_valid[1153]                      =   1'b0;
assign   tb_i_reset[1153]                      =   1'b0;
assign   tb_i_sop[1153]                        =   1'b0;
assign   tb_i_key_update[1153]                 =   1'b0;
assign   tb_i_key[1153]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1153]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1153]               =   1'b0;
assign   tb_i_rf_static_encrypt[1153]          =   1'b1;
assign   tb_i_clear_fault_flags[1153]          =   1'b0;
assign   tb_i_rf_static_aad_length[1153]       =   64'h0000000000000100;
assign   tb_i_aad[1153]                        =   tb_i_aad[1152];
assign   tb_i_rf_static_plaintext_length[1153] =   64'h0000000000000280;
assign   tb_i_plaintext[1153]                  =   tb_i_plaintext[1152];
assign   tb_o_valid[1153]                      =   1'b0;
assign   tb_o_sop[1153]                        =   1'b0;
assign   tb_o_ciphertext[1153]                 =   tb_o_ciphertext[1152];
assign   tb_o_tag_ready[1153]                  =   1'b0;
assign   tb_o_tag[1153]                        =   tb_o_tag[1152];

// CLK no. 1154/1240
// *************************************************
assign   tb_i_valid[1154]                      =   1'b0;
assign   tb_i_reset[1154]                      =   1'b0;
assign   tb_i_sop[1154]                        =   1'b0;
assign   tb_i_key_update[1154]                 =   1'b0;
assign   tb_i_key[1154]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1154]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1154]               =   1'b0;
assign   tb_i_rf_static_encrypt[1154]          =   1'b1;
assign   tb_i_clear_fault_flags[1154]          =   1'b0;
assign   tb_i_rf_static_aad_length[1154]       =   64'h0000000000000100;
assign   tb_i_aad[1154]                        =   tb_i_aad[1153];
assign   tb_i_rf_static_plaintext_length[1154] =   64'h0000000000000280;
assign   tb_i_plaintext[1154]                  =   tb_i_plaintext[1153];
assign   tb_o_valid[1154]                      =   1'b0;
assign   tb_o_sop[1154]                        =   1'b0;
assign   tb_o_ciphertext[1154]                 =   tb_o_ciphertext[1153];
assign   tb_o_tag_ready[1154]                  =   1'b0;
assign   tb_o_tag[1154]                        =   tb_o_tag[1153];

// CLK no. 1155/1240
// *************************************************
assign   tb_i_valid[1155]                      =   1'b0;
assign   tb_i_reset[1155]                      =   1'b0;
assign   tb_i_sop[1155]                        =   1'b0;
assign   tb_i_key_update[1155]                 =   1'b0;
assign   tb_i_key[1155]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1155]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1155]               =   1'b0;
assign   tb_i_rf_static_encrypt[1155]          =   1'b1;
assign   tb_i_clear_fault_flags[1155]          =   1'b0;
assign   tb_i_rf_static_aad_length[1155]       =   64'h0000000000000100;
assign   tb_i_aad[1155]                        =   tb_i_aad[1154];
assign   tb_i_rf_static_plaintext_length[1155] =   64'h0000000000000280;
assign   tb_i_plaintext[1155]                  =   tb_i_plaintext[1154];
assign   tb_o_valid[1155]                      =   1'b0;
assign   tb_o_sop[1155]                        =   1'b0;
assign   tb_o_ciphertext[1155]                 =   tb_o_ciphertext[1154];
assign   tb_o_tag_ready[1155]                  =   1'b0;
assign   tb_o_tag[1155]                        =   tb_o_tag[1154];

// CLK no. 1156/1240
// *************************************************
assign   tb_i_valid[1156]                      =   1'b0;
assign   tb_i_reset[1156]                      =   1'b0;
assign   tb_i_sop[1156]                        =   1'b0;
assign   tb_i_key_update[1156]                 =   1'b0;
assign   tb_i_key[1156]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1156]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1156]               =   1'b0;
assign   tb_i_rf_static_encrypt[1156]          =   1'b1;
assign   tb_i_clear_fault_flags[1156]          =   1'b0;
assign   tb_i_rf_static_aad_length[1156]       =   64'h0000000000000100;
assign   tb_i_aad[1156]                        =   tb_i_aad[1155];
assign   tb_i_rf_static_plaintext_length[1156] =   64'h0000000000000280;
assign   tb_i_plaintext[1156]                  =   tb_i_plaintext[1155];
assign   tb_o_valid[1156]                      =   1'b0;
assign   tb_o_sop[1156]                        =   1'b0;
assign   tb_o_ciphertext[1156]                 =   tb_o_ciphertext[1155];
assign   tb_o_tag_ready[1156]                  =   1'b0;
assign   tb_o_tag[1156]                        =   tb_o_tag[1155];

// CLK no. 1157/1240
// *************************************************
assign   tb_i_valid[1157]                      =   1'b0;
assign   tb_i_reset[1157]                      =   1'b0;
assign   tb_i_sop[1157]                        =   1'b0;
assign   tb_i_key_update[1157]                 =   1'b0;
assign   tb_i_key[1157]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1157]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1157]               =   1'b0;
assign   tb_i_rf_static_encrypt[1157]          =   1'b1;
assign   tb_i_clear_fault_flags[1157]          =   1'b0;
assign   tb_i_rf_static_aad_length[1157]       =   64'h0000000000000100;
assign   tb_i_aad[1157]                        =   tb_i_aad[1156];
assign   tb_i_rf_static_plaintext_length[1157] =   64'h0000000000000280;
assign   tb_i_plaintext[1157]                  =   tb_i_plaintext[1156];
assign   tb_o_valid[1157]                      =   1'b0;
assign   tb_o_sop[1157]                        =   1'b0;
assign   tb_o_ciphertext[1157]                 =   tb_o_ciphertext[1156];
assign   tb_o_tag_ready[1157]                  =   1'b0;
assign   tb_o_tag[1157]                        =   tb_o_tag[1156];

// CLK no. 1158/1240
// *************************************************
assign   tb_i_valid[1158]                      =   1'b0;
assign   tb_i_reset[1158]                      =   1'b0;
assign   tb_i_sop[1158]                        =   1'b0;
assign   tb_i_key_update[1158]                 =   1'b0;
assign   tb_i_key[1158]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1158]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1158]               =   1'b0;
assign   tb_i_rf_static_encrypt[1158]          =   1'b1;
assign   tb_i_clear_fault_flags[1158]          =   1'b0;
assign   tb_i_rf_static_aad_length[1158]       =   64'h0000000000000100;
assign   tb_i_aad[1158]                        =   tb_i_aad[1157];
assign   tb_i_rf_static_plaintext_length[1158] =   64'h0000000000000280;
assign   tb_i_plaintext[1158]                  =   tb_i_plaintext[1157];
assign   tb_o_valid[1158]                      =   1'b0;
assign   tb_o_sop[1158]                        =   1'b0;
assign   tb_o_ciphertext[1158]                 =   tb_o_ciphertext[1157];
assign   tb_o_tag_ready[1158]                  =   1'b0;
assign   tb_o_tag[1158]                        =   tb_o_tag[1157];

// CLK no. 1159/1240
// *************************************************
assign   tb_i_valid[1159]                      =   1'b0;
assign   tb_i_reset[1159]                      =   1'b0;
assign   tb_i_sop[1159]                        =   1'b0;
assign   tb_i_key_update[1159]                 =   1'b0;
assign   tb_i_key[1159]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1159]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1159]               =   1'b0;
assign   tb_i_rf_static_encrypt[1159]          =   1'b1;
assign   tb_i_clear_fault_flags[1159]          =   1'b0;
assign   tb_i_rf_static_aad_length[1159]       =   64'h0000000000000100;
assign   tb_i_aad[1159]                        =   tb_i_aad[1158];
assign   tb_i_rf_static_plaintext_length[1159] =   64'h0000000000000280;
assign   tb_i_plaintext[1159]                  =   tb_i_plaintext[1158];
assign   tb_o_valid[1159]                      =   1'b0;
assign   tb_o_sop[1159]                        =   1'b0;
assign   tb_o_ciphertext[1159]                 =   tb_o_ciphertext[1158];
assign   tb_o_tag_ready[1159]                  =   1'b0;
assign   tb_o_tag[1159]                        =   tb_o_tag[1158];

// CLK no. 1160/1240
// *************************************************
assign   tb_i_valid[1160]                      =   1'b0;
assign   tb_i_reset[1160]                      =   1'b0;
assign   tb_i_sop[1160]                        =   1'b0;
assign   tb_i_key_update[1160]                 =   1'b0;
assign   tb_i_key[1160]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1160]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1160]               =   1'b0;
assign   tb_i_rf_static_encrypt[1160]          =   1'b1;
assign   tb_i_clear_fault_flags[1160]          =   1'b0;
assign   tb_i_rf_static_aad_length[1160]       =   64'h0000000000000100;
assign   tb_i_aad[1160]                        =   tb_i_aad[1159];
assign   tb_i_rf_static_plaintext_length[1160] =   64'h0000000000000280;
assign   tb_i_plaintext[1160]                  =   tb_i_plaintext[1159];
assign   tb_o_valid[1160]                      =   1'b0;
assign   tb_o_sop[1160]                        =   1'b0;
assign   tb_o_ciphertext[1160]                 =   tb_o_ciphertext[1159];
assign   tb_o_tag_ready[1160]                  =   1'b0;
assign   tb_o_tag[1160]                        =   tb_o_tag[1159];

// CLK no. 1161/1240
// *************************************************
assign   tb_i_valid[1161]                      =   1'b0;
assign   tb_i_reset[1161]                      =   1'b0;
assign   tb_i_sop[1161]                        =   1'b0;
assign   tb_i_key_update[1161]                 =   1'b0;
assign   tb_i_key[1161]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1161]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1161]               =   1'b0;
assign   tb_i_rf_static_encrypt[1161]          =   1'b1;
assign   tb_i_clear_fault_flags[1161]          =   1'b0;
assign   tb_i_rf_static_aad_length[1161]       =   64'h0000000000000100;
assign   tb_i_aad[1161]                        =   tb_i_aad[1160];
assign   tb_i_rf_static_plaintext_length[1161] =   64'h0000000000000280;
assign   tb_i_plaintext[1161]                  =   tb_i_plaintext[1160];
assign   tb_o_valid[1161]                      =   1'b0;
assign   tb_o_sop[1161]                        =   1'b0;
assign   tb_o_ciphertext[1161]                 =   tb_o_ciphertext[1160];
assign   tb_o_tag_ready[1161]                  =   1'b0;
assign   tb_o_tag[1161]                        =   tb_o_tag[1160];

// CLK no. 1162/1240
// *************************************************
assign   tb_i_valid[1162]                      =   1'b0;
assign   tb_i_reset[1162]                      =   1'b0;
assign   tb_i_sop[1162]                        =   1'b0;
assign   tb_i_key_update[1162]                 =   1'b0;
assign   tb_i_key[1162]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1162]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1162]               =   1'b0;
assign   tb_i_rf_static_encrypt[1162]          =   1'b1;
assign   tb_i_clear_fault_flags[1162]          =   1'b0;
assign   tb_i_rf_static_aad_length[1162]       =   64'h0000000000000100;
assign   tb_i_aad[1162]                        =   tb_i_aad[1161];
assign   tb_i_rf_static_plaintext_length[1162] =   64'h0000000000000280;
assign   tb_i_plaintext[1162]                  =   tb_i_plaintext[1161];
assign   tb_o_valid[1162]                      =   1'b0;
assign   tb_o_sop[1162]                        =   1'b0;
assign   tb_o_ciphertext[1162]                 =   tb_o_ciphertext[1161];
assign   tb_o_tag_ready[1162]                  =   1'b0;
assign   tb_o_tag[1162]                        =   tb_o_tag[1161];

// CLK no. 1163/1240
// *************************************************
assign   tb_i_valid[1163]                      =   1'b0;
assign   tb_i_reset[1163]                      =   1'b0;
assign   tb_i_sop[1163]                        =   1'b0;
assign   tb_i_key_update[1163]                 =   1'b0;
assign   tb_i_key[1163]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1163]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1163]               =   1'b0;
assign   tb_i_rf_static_encrypt[1163]          =   1'b1;
assign   tb_i_clear_fault_flags[1163]          =   1'b0;
assign   tb_i_rf_static_aad_length[1163]       =   64'h0000000000000100;
assign   tb_i_aad[1163]                        =   tb_i_aad[1162];
assign   tb_i_rf_static_plaintext_length[1163] =   64'h0000000000000280;
assign   tb_i_plaintext[1163]                  =   tb_i_plaintext[1162];
assign   tb_o_valid[1163]                      =   1'b0;
assign   tb_o_sop[1163]                        =   1'b0;
assign   tb_o_ciphertext[1163]                 =   tb_o_ciphertext[1162];
assign   tb_o_tag_ready[1163]                  =   1'b0;
assign   tb_o_tag[1163]                        =   tb_o_tag[1162];

// CLK no. 1164/1240
// *************************************************
assign   tb_i_valid[1164]                      =   1'b0;
assign   tb_i_reset[1164]                      =   1'b0;
assign   tb_i_sop[1164]                        =   1'b0;
assign   tb_i_key_update[1164]                 =   1'b0;
assign   tb_i_key[1164]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1164]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1164]               =   1'b0;
assign   tb_i_rf_static_encrypt[1164]          =   1'b1;
assign   tb_i_clear_fault_flags[1164]          =   1'b0;
assign   tb_i_rf_static_aad_length[1164]       =   64'h0000000000000100;
assign   tb_i_aad[1164]                        =   tb_i_aad[1163];
assign   tb_i_rf_static_plaintext_length[1164] =   64'h0000000000000280;
assign   tb_i_plaintext[1164]                  =   tb_i_plaintext[1163];
assign   tb_o_valid[1164]                      =   1'b0;
assign   tb_o_sop[1164]                        =   1'b0;
assign   tb_o_ciphertext[1164]                 =   tb_o_ciphertext[1163];
assign   tb_o_tag_ready[1164]                  =   1'b0;
assign   tb_o_tag[1164]                        =   tb_o_tag[1163];

// CLK no. 1165/1240
// *************************************************
assign   tb_i_valid[1165]                      =   1'b0;
assign   tb_i_reset[1165]                      =   1'b0;
assign   tb_i_sop[1165]                        =   1'b0;
assign   tb_i_key_update[1165]                 =   1'b0;
assign   tb_i_key[1165]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1165]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1165]               =   1'b0;
assign   tb_i_rf_static_encrypt[1165]          =   1'b1;
assign   tb_i_clear_fault_flags[1165]          =   1'b0;
assign   tb_i_rf_static_aad_length[1165]       =   64'h0000000000000100;
assign   tb_i_aad[1165]                        =   tb_i_aad[1164];
assign   tb_i_rf_static_plaintext_length[1165] =   64'h0000000000000280;
assign   tb_i_plaintext[1165]                  =   tb_i_plaintext[1164];
assign   tb_o_valid[1165]                      =   1'b0;
assign   tb_o_sop[1165]                        =   1'b0;
assign   tb_o_ciphertext[1165]                 =   tb_o_ciphertext[1164];
assign   tb_o_tag_ready[1165]                  =   1'b0;
assign   tb_o_tag[1165]                        =   tb_o_tag[1164];

// CLK no. 1166/1240
// *************************************************
assign   tb_i_valid[1166]                      =   1'b0;
assign   tb_i_reset[1166]                      =   1'b0;
assign   tb_i_sop[1166]                        =   1'b0;
assign   tb_i_key_update[1166]                 =   1'b0;
assign   tb_i_key[1166]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1166]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1166]               =   1'b0;
assign   tb_i_rf_static_encrypt[1166]          =   1'b1;
assign   tb_i_clear_fault_flags[1166]          =   1'b0;
assign   tb_i_rf_static_aad_length[1166]       =   64'h0000000000000100;
assign   tb_i_aad[1166]                        =   tb_i_aad[1165];
assign   tb_i_rf_static_plaintext_length[1166] =   64'h0000000000000280;
assign   tb_i_plaintext[1166]                  =   tb_i_plaintext[1165];
assign   tb_o_valid[1166]                      =   1'b0;
assign   tb_o_sop[1166]                        =   1'b0;
assign   tb_o_ciphertext[1166]                 =   tb_o_ciphertext[1165];
assign   tb_o_tag_ready[1166]                  =   1'b0;
assign   tb_o_tag[1166]                        =   tb_o_tag[1165];

// CLK no. 1167/1240
// *************************************************
assign   tb_i_valid[1167]                      =   1'b0;
assign   tb_i_reset[1167]                      =   1'b0;
assign   tb_i_sop[1167]                        =   1'b0;
assign   tb_i_key_update[1167]                 =   1'b0;
assign   tb_i_key[1167]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1167]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1167]               =   1'b0;
assign   tb_i_rf_static_encrypt[1167]          =   1'b1;
assign   tb_i_clear_fault_flags[1167]          =   1'b0;
assign   tb_i_rf_static_aad_length[1167]       =   64'h0000000000000100;
assign   tb_i_aad[1167]                        =   tb_i_aad[1166];
assign   tb_i_rf_static_plaintext_length[1167] =   64'h0000000000000280;
assign   tb_i_plaintext[1167]                  =   tb_i_plaintext[1166];
assign   tb_o_valid[1167]                      =   1'b0;
assign   tb_o_sop[1167]                        =   1'b0;
assign   tb_o_ciphertext[1167]                 =   tb_o_ciphertext[1166];
assign   tb_o_tag_ready[1167]                  =   1'b0;
assign   tb_o_tag[1167]                        =   tb_o_tag[1166];

// CLK no. 1168/1240
// *************************************************
assign   tb_i_valid[1168]                      =   1'b0;
assign   tb_i_reset[1168]                      =   1'b0;
assign   tb_i_sop[1168]                        =   1'b0;
assign   tb_i_key_update[1168]                 =   1'b0;
assign   tb_i_key[1168]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1168]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1168]               =   1'b0;
assign   tb_i_rf_static_encrypt[1168]          =   1'b1;
assign   tb_i_clear_fault_flags[1168]          =   1'b0;
assign   tb_i_rf_static_aad_length[1168]       =   64'h0000000000000100;
assign   tb_i_aad[1168]                        =   tb_i_aad[1167];
assign   tb_i_rf_static_plaintext_length[1168] =   64'h0000000000000280;
assign   tb_i_plaintext[1168]                  =   tb_i_plaintext[1167];
assign   tb_o_valid[1168]                      =   1'b1;
assign   tb_o_sop[1168]                        =   1'b1;
assign   tb_o_ciphertext[1168]                 =   256'h462cd4d4b6fc29e7e32514b55d3f512b2e4fa72ae0ff2a311ea9936a4c47d4af;
assign   tb_o_tag_ready[1168]                  =   1'b0;
assign   tb_o_tag[1168]                        =   tb_o_tag[1167];

// CLK no. 1169/1240
// *************************************************
assign   tb_i_valid[1169]                      =   1'b0;
assign   tb_i_reset[1169]                      =   1'b0;
assign   tb_i_sop[1169]                        =   1'b0;
assign   tb_i_key_update[1169]                 =   1'b0;
assign   tb_i_key[1169]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1169]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1169]               =   1'b0;
assign   tb_i_rf_static_encrypt[1169]          =   1'b1;
assign   tb_i_clear_fault_flags[1169]          =   1'b0;
assign   tb_i_rf_static_aad_length[1169]       =   64'h0000000000000100;
assign   tb_i_aad[1169]                        =   tb_i_aad[1168];
assign   tb_i_rf_static_plaintext_length[1169] =   64'h0000000000000280;
assign   tb_i_plaintext[1169]                  =   tb_i_plaintext[1168];
assign   tb_o_valid[1169]                      =   1'b1;
assign   tb_o_sop[1169]                        =   1'b0;
assign   tb_o_ciphertext[1169]                 =   256'h04c54e92631864a248520fbc0b5c6ba030ed4e229f26b508c6a0dc111d868535;
assign   tb_o_tag_ready[1169]                  =   1'b0;
assign   tb_o_tag[1169]                        =   tb_o_tag[1168];

// CLK no. 1170/1240
// *************************************************
assign   tb_i_valid[1170]                      =   1'b0;
assign   tb_i_reset[1170]                      =   1'b0;
assign   tb_i_sop[1170]                        =   1'b0;
assign   tb_i_key_update[1170]                 =   1'b0;
assign   tb_i_key[1170]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1170]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1170]               =   1'b0;
assign   tb_i_rf_static_encrypt[1170]          =   1'b1;
assign   tb_i_clear_fault_flags[1170]          =   1'b0;
assign   tb_i_rf_static_aad_length[1170]       =   64'h0000000000000100;
assign   tb_i_aad[1170]                        =   tb_i_aad[1169];
assign   tb_i_rf_static_plaintext_length[1170] =   64'h0000000000000280;
assign   tb_i_plaintext[1170]                  =   tb_i_plaintext[1169];
assign   tb_o_valid[1170]                      =   1'b1;
assign   tb_o_sop[1170]                        =   1'b0;
assign   tb_o_ciphertext[1170]                 =   256'h923c53664e92bde609303ba103309de7;
assign   tb_o_tag_ready[1170]                  =   1'b0;
assign   tb_o_tag[1170]                        =   tb_o_tag[1169];

// CLK no. 1171/1240
// *************************************************
assign   tb_i_valid[1171]                      =   1'b0;
assign   tb_i_reset[1171]                      =   1'b0;
assign   tb_i_sop[1171]                        =   1'b0;
assign   tb_i_key_update[1171]                 =   1'b0;
assign   tb_i_key[1171]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1171]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1171]               =   1'b0;
assign   tb_i_rf_static_encrypt[1171]          =   1'b1;
assign   tb_i_clear_fault_flags[1171]          =   1'b0;
assign   tb_i_rf_static_aad_length[1171]       =   64'h0000000000000100;
assign   tb_i_aad[1171]                        =   tb_i_aad[1170];
assign   tb_i_rf_static_plaintext_length[1171] =   64'h0000000000000280;
assign   tb_i_plaintext[1171]                  =   tb_i_plaintext[1170];
assign   tb_o_valid[1171]                      =   1'b0;
assign   tb_o_sop[1171]                        =   1'b0;
assign   tb_o_ciphertext[1171]                 =   tb_o_ciphertext[1170];
assign   tb_o_tag_ready[1171]                  =   1'b0;
assign   tb_o_tag[1171]                        =   tb_o_tag[1170];

// CLK no. 1172/1240
// *************************************************
assign   tb_i_valid[1172]                      =   1'b0;
assign   tb_i_reset[1172]                      =   1'b0;
assign   tb_i_sop[1172]                        =   1'b0;
assign   tb_i_key_update[1172]                 =   1'b0;
assign   tb_i_key[1172]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1172]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1172]               =   1'b0;
assign   tb_i_rf_static_encrypt[1172]          =   1'b1;
assign   tb_i_clear_fault_flags[1172]          =   1'b0;
assign   tb_i_rf_static_aad_length[1172]       =   64'h0000000000000100;
assign   tb_i_aad[1172]                        =   tb_i_aad[1171];
assign   tb_i_rf_static_plaintext_length[1172] =   64'h0000000000000280;
assign   tb_i_plaintext[1172]                  =   tb_i_plaintext[1171];
assign   tb_o_valid[1172]                      =   1'b0;
assign   tb_o_sop[1172]                        =   1'b0;
assign   tb_o_ciphertext[1172]                 =   tb_o_ciphertext[1171];
assign   tb_o_tag_ready[1172]                  =   1'b0;
assign   tb_o_tag[1172]                        =   tb_o_tag[1171];

// CLK no. 1173/1240
// *************************************************
assign   tb_i_valid[1173]                      =   1'b0;
assign   tb_i_reset[1173]                      =   1'b0;
assign   tb_i_sop[1173]                        =   1'b0;
assign   tb_i_key_update[1173]                 =   1'b0;
assign   tb_i_key[1173]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1173]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1173]               =   1'b0;
assign   tb_i_rf_static_encrypt[1173]          =   1'b1;
assign   tb_i_clear_fault_flags[1173]          =   1'b0;
assign   tb_i_rf_static_aad_length[1173]       =   64'h0000000000000100;
assign   tb_i_aad[1173]                        =   tb_i_aad[1172];
assign   tb_i_rf_static_plaintext_length[1173] =   64'h0000000000000280;
assign   tb_i_plaintext[1173]                  =   tb_i_plaintext[1172];
assign   tb_o_valid[1173]                      =   1'b0;
assign   tb_o_sop[1173]                        =   1'b0;
assign   tb_o_ciphertext[1173]                 =   tb_o_ciphertext[1172];
assign   tb_o_tag_ready[1173]                  =   1'b0;
assign   tb_o_tag[1173]                        =   tb_o_tag[1172];

// CLK no. 1174/1240
// *************************************************
assign   tb_i_valid[1174]                      =   1'b0;
assign   tb_i_reset[1174]                      =   1'b0;
assign   tb_i_sop[1174]                        =   1'b0;
assign   tb_i_key_update[1174]                 =   1'b0;
assign   tb_i_key[1174]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1174]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1174]               =   1'b0;
assign   tb_i_rf_static_encrypt[1174]          =   1'b1;
assign   tb_i_clear_fault_flags[1174]          =   1'b0;
assign   tb_i_rf_static_aad_length[1174]       =   64'h0000000000000100;
assign   tb_i_aad[1174]                        =   tb_i_aad[1173];
assign   tb_i_rf_static_plaintext_length[1174] =   64'h0000000000000280;
assign   tb_i_plaintext[1174]                  =   tb_i_plaintext[1173];
assign   tb_o_valid[1174]                      =   1'b0;
assign   tb_o_sop[1174]                        =   1'b0;
assign   tb_o_ciphertext[1174]                 =   tb_o_ciphertext[1173];
assign   tb_o_tag_ready[1174]                  =   1'b0;
assign   tb_o_tag[1174]                        =   tb_o_tag[1173];

// CLK no. 1175/1240
// *************************************************
assign   tb_i_valid[1175]                      =   1'b0;
assign   tb_i_reset[1175]                      =   1'b0;
assign   tb_i_sop[1175]                        =   1'b0;
assign   tb_i_key_update[1175]                 =   1'b0;
assign   tb_i_key[1175]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1175]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1175]               =   1'b0;
assign   tb_i_rf_static_encrypt[1175]          =   1'b1;
assign   tb_i_clear_fault_flags[1175]          =   1'b0;
assign   tb_i_rf_static_aad_length[1175]       =   64'h0000000000000100;
assign   tb_i_aad[1175]                        =   tb_i_aad[1174];
assign   tb_i_rf_static_plaintext_length[1175] =   64'h0000000000000280;
assign   tb_i_plaintext[1175]                  =   tb_i_plaintext[1174];
assign   tb_o_valid[1175]                      =   1'b0;
assign   tb_o_sop[1175]                        =   1'b0;
assign   tb_o_ciphertext[1175]                 =   tb_o_ciphertext[1174];
assign   tb_o_tag_ready[1175]                  =   1'b0;
assign   tb_o_tag[1175]                        =   tb_o_tag[1174];

// CLK no. 1176/1240
// *************************************************
assign   tb_i_valid[1176]                      =   1'b0;
assign   tb_i_reset[1176]                      =   1'b0;
assign   tb_i_sop[1176]                        =   1'b0;
assign   tb_i_key_update[1176]                 =   1'b0;
assign   tb_i_key[1176]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1176]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1176]               =   1'b0;
assign   tb_i_rf_static_encrypt[1176]          =   1'b1;
assign   tb_i_clear_fault_flags[1176]          =   1'b0;
assign   tb_i_rf_static_aad_length[1176]       =   64'h0000000000000100;
assign   tb_i_aad[1176]                        =   tb_i_aad[1175];
assign   tb_i_rf_static_plaintext_length[1176] =   64'h0000000000000280;
assign   tb_i_plaintext[1176]                  =   tb_i_plaintext[1175];
assign   tb_o_valid[1176]                      =   1'b0;
assign   tb_o_sop[1176]                        =   1'b0;
assign   tb_o_ciphertext[1176]                 =   tb_o_ciphertext[1175];
assign   tb_o_tag_ready[1176]                  =   1'b0;
assign   tb_o_tag[1176]                        =   tb_o_tag[1175];

// CLK no. 1177/1240
// *************************************************
assign   tb_i_valid[1177]                      =   1'b0;
assign   tb_i_reset[1177]                      =   1'b0;
assign   tb_i_sop[1177]                        =   1'b0;
assign   tb_i_key_update[1177]                 =   1'b0;
assign   tb_i_key[1177]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1177]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1177]               =   1'b0;
assign   tb_i_rf_static_encrypt[1177]          =   1'b1;
assign   tb_i_clear_fault_flags[1177]          =   1'b0;
assign   tb_i_rf_static_aad_length[1177]       =   64'h0000000000000100;
assign   tb_i_aad[1177]                        =   tb_i_aad[1176];
assign   tb_i_rf_static_plaintext_length[1177] =   64'h0000000000000280;
assign   tb_i_plaintext[1177]                  =   tb_i_plaintext[1176];
assign   tb_o_valid[1177]                      =   1'b0;
assign   tb_o_sop[1177]                        =   1'b0;
assign   tb_o_ciphertext[1177]                 =   tb_o_ciphertext[1176];
assign   tb_o_tag_ready[1177]                  =   1'b0;
assign   tb_o_tag[1177]                        =   tb_o_tag[1176];

// CLK no. 1178/1240
// *************************************************
assign   tb_i_valid[1178]                      =   1'b0;
assign   tb_i_reset[1178]                      =   1'b0;
assign   tb_i_sop[1178]                        =   1'b0;
assign   tb_i_key_update[1178]                 =   1'b0;
assign   tb_i_key[1178]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1178]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1178]               =   1'b0;
assign   tb_i_rf_static_encrypt[1178]          =   1'b1;
assign   tb_i_clear_fault_flags[1178]          =   1'b0;
assign   tb_i_rf_static_aad_length[1178]       =   64'h0000000000000100;
assign   tb_i_aad[1178]                        =   tb_i_aad[1177];
assign   tb_i_rf_static_plaintext_length[1178] =   64'h0000000000000280;
assign   tb_i_plaintext[1178]                  =   tb_i_plaintext[1177];
assign   tb_o_valid[1178]                      =   1'b0;
assign   tb_o_sop[1178]                        =   1'b0;
assign   tb_o_ciphertext[1178]                 =   tb_o_ciphertext[1177];
assign   tb_o_tag_ready[1178]                  =   1'b1;
assign   tb_o_tag[1178]                        =   128'hd8f2fe9f17e3b1ca6cb67951bb4e37c7;

// CLK no. 1179/1240
// *************************************************
assign   tb_i_valid[1179]                      =   1'b0;
assign   tb_i_reset[1179]                      =   1'b0;
assign   tb_i_sop[1179]                        =   1'b0;
assign   tb_i_key_update[1179]                 =   1'b0;
assign   tb_i_key[1179]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1179]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1179]               =   1'b0;
assign   tb_i_rf_static_encrypt[1179]          =   1'b1;
assign   tb_i_clear_fault_flags[1179]          =   1'b0;
assign   tb_i_rf_static_aad_length[1179]       =   64'h0000000000000100;
assign   tb_i_aad[1179]                        =   tb_i_aad[1178];
assign   tb_i_rf_static_plaintext_length[1179] =   64'h0000000000000280;
assign   tb_i_plaintext[1179]                  =   tb_i_plaintext[1178];
assign   tb_o_valid[1179]                      =   1'b0;
assign   tb_o_sop[1179]                        =   1'b0;
assign   tb_o_ciphertext[1179]                 =   tb_o_ciphertext[1178];
assign   tb_o_tag_ready[1179]                  =   1'b0;
assign   tb_o_tag[1179]                        =   tb_o_tag[1178];

// CLK no. 1180/1240
// *************************************************
assign   tb_i_valid[1180]                      =   1'b0;
assign   tb_i_reset[1180]                      =   1'b0;
assign   tb_i_sop[1180]                        =   1'b0;
assign   tb_i_key_update[1180]                 =   1'b0;
assign   tb_i_key[1180]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1180]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1180]               =   1'b0;
assign   tb_i_rf_static_encrypt[1180]          =   1'b1;
assign   tb_i_clear_fault_flags[1180]          =   1'b0;
assign   tb_i_rf_static_aad_length[1180]       =   64'h0000000000000100;
assign   tb_i_aad[1180]                        =   tb_i_aad[1179];
assign   tb_i_rf_static_plaintext_length[1180] =   64'h0000000000000280;
assign   tb_i_plaintext[1180]                  =   tb_i_plaintext[1179];
assign   tb_o_valid[1180]                      =   1'b0;
assign   tb_o_sop[1180]                        =   1'b0;
assign   tb_o_ciphertext[1180]                 =   tb_o_ciphertext[1179];
assign   tb_o_tag_ready[1180]                  =   1'b0;
assign   tb_o_tag[1180]                        =   tb_o_tag[1179];

// CLK no. 1181/1240
// *************************************************
assign   tb_i_valid[1181]                      =   1'b0;
assign   tb_i_reset[1181]                      =   1'b0;
assign   tb_i_sop[1181]                        =   1'b1;
assign   tb_i_key_update[1181]                 =   1'b0;
assign   tb_i_key[1181]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1181]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1181]               =   1'b0;
assign   tb_i_rf_static_encrypt[1181]          =   1'b1;
assign   tb_i_clear_fault_flags[1181]          =   1'b0;
assign   tb_i_rf_static_aad_length[1181]       =   64'h0000000000000100;
assign   tb_i_aad[1181]                        =   tb_i_aad[1180];
assign   tb_i_rf_static_plaintext_length[1181] =   64'h0000000000000280;
assign   tb_i_plaintext[1181]                  =   tb_i_plaintext[1180];
assign   tb_o_valid[1181]                      =   1'b0;
assign   tb_o_sop[1181]                        =   1'b0;
assign   tb_o_ciphertext[1181]                 =   tb_o_ciphertext[1180];
assign   tb_o_tag_ready[1181]                  =   1'b0;
assign   tb_o_tag[1181]                        =   tb_o_tag[1180];

// CLK no. 1182/1240
// *************************************************
assign   tb_i_valid[1182]                      =   1'b1;
assign   tb_i_reset[1182]                      =   1'b0;
assign   tb_i_sop[1182]                        =   1'b0;
assign   tb_i_key_update[1182]                 =   1'b0;
assign   tb_i_key[1182]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1182]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1182]               =   1'b0;
assign   tb_i_rf_static_encrypt[1182]          =   1'b1;
assign   tb_i_clear_fault_flags[1182]          =   1'b0;
assign   tb_i_rf_static_aad_length[1182]       =   64'h0000000000000100;
assign   tb_i_aad[1182]                        =   256'h31e6772f05039bf89afe4858e13a0866700d6b8e13fadf582e31b6b9431232cc;
assign   tb_i_rf_static_plaintext_length[1182] =   64'h0000000000000280;
assign   tb_i_plaintext[1182]                  =   tb_i_plaintext[1181];
assign   tb_o_valid[1182]                      =   1'b0;
assign   tb_o_sop[1182]                        =   1'b0;
assign   tb_o_ciphertext[1182]                 =   tb_o_ciphertext[1181];
assign   tb_o_tag_ready[1182]                  =   1'b0;
assign   tb_o_tag[1182]                        =   tb_o_tag[1181];

// CLK no. 1183/1240
// *************************************************
assign   tb_i_valid[1183]                      =   1'b1;
assign   tb_i_reset[1183]                      =   1'b0;
assign   tb_i_sop[1183]                        =   1'b0;
assign   tb_i_key_update[1183]                 =   1'b0;
assign   tb_i_key[1183]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1183]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1183]               =   1'b0;
assign   tb_i_rf_static_encrypt[1183]          =   1'b1;
assign   tb_i_clear_fault_flags[1183]          =   1'b0;
assign   tb_i_rf_static_aad_length[1183]       =   64'h0000000000000100;
assign   tb_i_aad[1183]                        =   tb_i_aad[1182];
assign   tb_i_rf_static_plaintext_length[1183] =   64'h0000000000000280;
assign   tb_i_plaintext[1183]                  =   256'h4caac8ca7c16a243c66f263d43f930ab81f7eae24596038e09bb89f750b916a5;
assign   tb_o_valid[1183]                      =   1'b0;
assign   tb_o_sop[1183]                        =   1'b0;
assign   tb_o_ciphertext[1183]                 =   tb_o_ciphertext[1182];
assign   tb_o_tag_ready[1183]                  =   1'b0;
assign   tb_o_tag[1183]                        =   tb_o_tag[1182];

// CLK no. 1184/1240
// *************************************************
assign   tb_i_valid[1184]                      =   1'b1;
assign   tb_i_reset[1184]                      =   1'b0;
assign   tb_i_sop[1184]                        =   1'b0;
assign   tb_i_key_update[1184]                 =   1'b0;
assign   tb_i_key[1184]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1184]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1184]               =   1'b0;
assign   tb_i_rf_static_encrypt[1184]          =   1'b1;
assign   tb_i_clear_fault_flags[1184]          =   1'b0;
assign   tb_i_rf_static_aad_length[1184]       =   64'h0000000000000100;
assign   tb_i_aad[1184]                        =   tb_i_aad[1183];
assign   tb_i_rf_static_plaintext_length[1184] =   64'h0000000000000280;
assign   tb_i_plaintext[1184]                  =   256'hefd6a67631a9f96f4d3e9d7c4ad352d87d390cb9654d0a281ce6ff13602c9380;
assign   tb_o_valid[1184]                      =   1'b0;
assign   tb_o_sop[1184]                        =   1'b0;
assign   tb_o_ciphertext[1184]                 =   tb_o_ciphertext[1183];
assign   tb_o_tag_ready[1184]                  =   1'b0;
assign   tb_o_tag[1184]                        =   tb_o_tag[1183];

// CLK no. 1185/1240
// *************************************************
assign   tb_i_valid[1185]                      =   1'b1;
assign   tb_i_reset[1185]                      =   1'b0;
assign   tb_i_sop[1185]                        =   1'b0;
assign   tb_i_key_update[1185]                 =   1'b0;
assign   tb_i_key[1185]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1185]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1185]               =   1'b0;
assign   tb_i_rf_static_encrypt[1185]          =   1'b1;
assign   tb_i_clear_fault_flags[1185]          =   1'b0;
assign   tb_i_rf_static_aad_length[1185]       =   64'h0000000000000100;
assign   tb_i_aad[1185]                        =   tb_i_aad[1184];
assign   tb_i_rf_static_plaintext_length[1185] =   64'h0000000000000280;
assign   tb_i_plaintext[1185]                  =   256'h578271150975701168055e37a262ca56;
assign   tb_o_valid[1185]                      =   1'b0;
assign   tb_o_sop[1185]                        =   1'b0;
assign   tb_o_ciphertext[1185]                 =   tb_o_ciphertext[1184];
assign   tb_o_tag_ready[1185]                  =   1'b0;
assign   tb_o_tag[1185]                        =   tb_o_tag[1184];

// CLK no. 1186/1240
// *************************************************
assign   tb_i_valid[1186]                      =   1'b0;
assign   tb_i_reset[1186]                      =   1'b0;
assign   tb_i_sop[1186]                        =   1'b0;
assign   tb_i_key_update[1186]                 =   1'b0;
assign   tb_i_key[1186]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1186]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1186]               =   1'b0;
assign   tb_i_rf_static_encrypt[1186]          =   1'b1;
assign   tb_i_clear_fault_flags[1186]          =   1'b0;
assign   tb_i_rf_static_aad_length[1186]       =   64'h0000000000000100;
assign   tb_i_aad[1186]                        =   tb_i_aad[1185];
assign   tb_i_rf_static_plaintext_length[1186] =   64'h0000000000000280;
assign   tb_i_plaintext[1186]                  =   tb_i_plaintext[1185];
assign   tb_o_valid[1186]                      =   1'b0;
assign   tb_o_sop[1186]                        =   1'b0;
assign   tb_o_ciphertext[1186]                 =   tb_o_ciphertext[1185];
assign   tb_o_tag_ready[1186]                  =   1'b0;
assign   tb_o_tag[1186]                        =   tb_o_tag[1185];

// CLK no. 1187/1240
// *************************************************
assign   tb_i_valid[1187]                      =   1'b0;
assign   tb_i_reset[1187]                      =   1'b0;
assign   tb_i_sop[1187]                        =   1'b0;
assign   tb_i_key_update[1187]                 =   1'b0;
assign   tb_i_key[1187]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1187]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1187]               =   1'b0;
assign   tb_i_rf_static_encrypt[1187]          =   1'b1;
assign   tb_i_clear_fault_flags[1187]          =   1'b0;
assign   tb_i_rf_static_aad_length[1187]       =   64'h0000000000000100;
assign   tb_i_aad[1187]                        =   tb_i_aad[1186];
assign   tb_i_rf_static_plaintext_length[1187] =   64'h0000000000000280;
assign   tb_i_plaintext[1187]                  =   tb_i_plaintext[1186];
assign   tb_o_valid[1187]                      =   1'b0;
assign   tb_o_sop[1187]                        =   1'b0;
assign   tb_o_ciphertext[1187]                 =   tb_o_ciphertext[1186];
assign   tb_o_tag_ready[1187]                  =   1'b0;
assign   tb_o_tag[1187]                        =   tb_o_tag[1186];

// CLK no. 1188/1240
// *************************************************
assign   tb_i_valid[1188]                      =   1'b0;
assign   tb_i_reset[1188]                      =   1'b0;
assign   tb_i_sop[1188]                        =   1'b0;
assign   tb_i_key_update[1188]                 =   1'b0;
assign   tb_i_key[1188]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1188]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1188]               =   1'b0;
assign   tb_i_rf_static_encrypt[1188]          =   1'b1;
assign   tb_i_clear_fault_flags[1188]          =   1'b0;
assign   tb_i_rf_static_aad_length[1188]       =   64'h0000000000000100;
assign   tb_i_aad[1188]                        =   tb_i_aad[1187];
assign   tb_i_rf_static_plaintext_length[1188] =   64'h0000000000000280;
assign   tb_i_plaintext[1188]                  =   tb_i_plaintext[1187];
assign   tb_o_valid[1188]                      =   1'b0;
assign   tb_o_sop[1188]                        =   1'b0;
assign   tb_o_ciphertext[1188]                 =   tb_o_ciphertext[1187];
assign   tb_o_tag_ready[1188]                  =   1'b0;
assign   tb_o_tag[1188]                        =   tb_o_tag[1187];

// CLK no. 1189/1240
// *************************************************
assign   tb_i_valid[1189]                      =   1'b0;
assign   tb_i_reset[1189]                      =   1'b0;
assign   tb_i_sop[1189]                        =   1'b0;
assign   tb_i_key_update[1189]                 =   1'b0;
assign   tb_i_key[1189]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1189]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1189]               =   1'b0;
assign   tb_i_rf_static_encrypt[1189]          =   1'b1;
assign   tb_i_clear_fault_flags[1189]          =   1'b0;
assign   tb_i_rf_static_aad_length[1189]       =   64'h0000000000000100;
assign   tb_i_aad[1189]                        =   tb_i_aad[1188];
assign   tb_i_rf_static_plaintext_length[1189] =   64'h0000000000000280;
assign   tb_i_plaintext[1189]                  =   tb_i_plaintext[1188];
assign   tb_o_valid[1189]                      =   1'b0;
assign   tb_o_sop[1189]                        =   1'b0;
assign   tb_o_ciphertext[1189]                 =   tb_o_ciphertext[1188];
assign   tb_o_tag_ready[1189]                  =   1'b0;
assign   tb_o_tag[1189]                        =   tb_o_tag[1188];

// CLK no. 1190/1240
// *************************************************
assign   tb_i_valid[1190]                      =   1'b0;
assign   tb_i_reset[1190]                      =   1'b0;
assign   tb_i_sop[1190]                        =   1'b0;
assign   tb_i_key_update[1190]                 =   1'b0;
assign   tb_i_key[1190]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1190]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1190]               =   1'b0;
assign   tb_i_rf_static_encrypt[1190]          =   1'b1;
assign   tb_i_clear_fault_flags[1190]          =   1'b0;
assign   tb_i_rf_static_aad_length[1190]       =   64'h0000000000000100;
assign   tb_i_aad[1190]                        =   tb_i_aad[1189];
assign   tb_i_rf_static_plaintext_length[1190] =   64'h0000000000000280;
assign   tb_i_plaintext[1190]                  =   tb_i_plaintext[1189];
assign   tb_o_valid[1190]                      =   1'b0;
assign   tb_o_sop[1190]                        =   1'b0;
assign   tb_o_ciphertext[1190]                 =   tb_o_ciphertext[1189];
assign   tb_o_tag_ready[1190]                  =   1'b0;
assign   tb_o_tag[1190]                        =   tb_o_tag[1189];

// CLK no. 1191/1240
// *************************************************
assign   tb_i_valid[1191]                      =   1'b0;
assign   tb_i_reset[1191]                      =   1'b0;
assign   tb_i_sop[1191]                        =   1'b0;
assign   tb_i_key_update[1191]                 =   1'b0;
assign   tb_i_key[1191]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1191]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1191]               =   1'b0;
assign   tb_i_rf_static_encrypt[1191]          =   1'b1;
assign   tb_i_clear_fault_flags[1191]          =   1'b0;
assign   tb_i_rf_static_aad_length[1191]       =   64'h0000000000000100;
assign   tb_i_aad[1191]                        =   tb_i_aad[1190];
assign   tb_i_rf_static_plaintext_length[1191] =   64'h0000000000000280;
assign   tb_i_plaintext[1191]                  =   tb_i_plaintext[1190];
assign   tb_o_valid[1191]                      =   1'b0;
assign   tb_o_sop[1191]                        =   1'b0;
assign   tb_o_ciphertext[1191]                 =   tb_o_ciphertext[1190];
assign   tb_o_tag_ready[1191]                  =   1'b0;
assign   tb_o_tag[1191]                        =   tb_o_tag[1190];

// CLK no. 1192/1240
// *************************************************
assign   tb_i_valid[1192]                      =   1'b0;
assign   tb_i_reset[1192]                      =   1'b0;
assign   tb_i_sop[1192]                        =   1'b0;
assign   tb_i_key_update[1192]                 =   1'b0;
assign   tb_i_key[1192]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1192]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1192]               =   1'b0;
assign   tb_i_rf_static_encrypt[1192]          =   1'b1;
assign   tb_i_clear_fault_flags[1192]          =   1'b0;
assign   tb_i_rf_static_aad_length[1192]       =   64'h0000000000000100;
assign   tb_i_aad[1192]                        =   tb_i_aad[1191];
assign   tb_i_rf_static_plaintext_length[1192] =   64'h0000000000000280;
assign   tb_i_plaintext[1192]                  =   tb_i_plaintext[1191];
assign   tb_o_valid[1192]                      =   1'b0;
assign   tb_o_sop[1192]                        =   1'b0;
assign   tb_o_ciphertext[1192]                 =   tb_o_ciphertext[1191];
assign   tb_o_tag_ready[1192]                  =   1'b0;
assign   tb_o_tag[1192]                        =   tb_o_tag[1191];

// CLK no. 1193/1240
// *************************************************
assign   tb_i_valid[1193]                      =   1'b0;
assign   tb_i_reset[1193]                      =   1'b0;
assign   tb_i_sop[1193]                        =   1'b0;
assign   tb_i_key_update[1193]                 =   1'b0;
assign   tb_i_key[1193]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1193]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1193]               =   1'b0;
assign   tb_i_rf_static_encrypt[1193]          =   1'b1;
assign   tb_i_clear_fault_flags[1193]          =   1'b0;
assign   tb_i_rf_static_aad_length[1193]       =   64'h0000000000000100;
assign   tb_i_aad[1193]                        =   tb_i_aad[1192];
assign   tb_i_rf_static_plaintext_length[1193] =   64'h0000000000000280;
assign   tb_i_plaintext[1193]                  =   tb_i_plaintext[1192];
assign   tb_o_valid[1193]                      =   1'b0;
assign   tb_o_sop[1193]                        =   1'b0;
assign   tb_o_ciphertext[1193]                 =   tb_o_ciphertext[1192];
assign   tb_o_tag_ready[1193]                  =   1'b0;
assign   tb_o_tag[1193]                        =   tb_o_tag[1192];

// CLK no. 1194/1240
// *************************************************
assign   tb_i_valid[1194]                      =   1'b0;
assign   tb_i_reset[1194]                      =   1'b0;
assign   tb_i_sop[1194]                        =   1'b0;
assign   tb_i_key_update[1194]                 =   1'b0;
assign   tb_i_key[1194]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1194]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1194]               =   1'b0;
assign   tb_i_rf_static_encrypt[1194]          =   1'b1;
assign   tb_i_clear_fault_flags[1194]          =   1'b0;
assign   tb_i_rf_static_aad_length[1194]       =   64'h0000000000000100;
assign   tb_i_aad[1194]                        =   tb_i_aad[1193];
assign   tb_i_rf_static_plaintext_length[1194] =   64'h0000000000000280;
assign   tb_i_plaintext[1194]                  =   tb_i_plaintext[1193];
assign   tb_o_valid[1194]                      =   1'b0;
assign   tb_o_sop[1194]                        =   1'b0;
assign   tb_o_ciphertext[1194]                 =   tb_o_ciphertext[1193];
assign   tb_o_tag_ready[1194]                  =   1'b0;
assign   tb_o_tag[1194]                        =   tb_o_tag[1193];

// CLK no. 1195/1240
// *************************************************
assign   tb_i_valid[1195]                      =   1'b0;
assign   tb_i_reset[1195]                      =   1'b0;
assign   tb_i_sop[1195]                        =   1'b0;
assign   tb_i_key_update[1195]                 =   1'b0;
assign   tb_i_key[1195]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1195]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1195]               =   1'b0;
assign   tb_i_rf_static_encrypt[1195]          =   1'b1;
assign   tb_i_clear_fault_flags[1195]          =   1'b0;
assign   tb_i_rf_static_aad_length[1195]       =   64'h0000000000000100;
assign   tb_i_aad[1195]                        =   tb_i_aad[1194];
assign   tb_i_rf_static_plaintext_length[1195] =   64'h0000000000000280;
assign   tb_i_plaintext[1195]                  =   tb_i_plaintext[1194];
assign   tb_o_valid[1195]                      =   1'b0;
assign   tb_o_sop[1195]                        =   1'b0;
assign   tb_o_ciphertext[1195]                 =   tb_o_ciphertext[1194];
assign   tb_o_tag_ready[1195]                  =   1'b0;
assign   tb_o_tag[1195]                        =   tb_o_tag[1194];

// CLK no. 1196/1240
// *************************************************
assign   tb_i_valid[1196]                      =   1'b0;
assign   tb_i_reset[1196]                      =   1'b0;
assign   tb_i_sop[1196]                        =   1'b0;
assign   tb_i_key_update[1196]                 =   1'b0;
assign   tb_i_key[1196]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1196]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1196]               =   1'b0;
assign   tb_i_rf_static_encrypt[1196]          =   1'b1;
assign   tb_i_clear_fault_flags[1196]          =   1'b0;
assign   tb_i_rf_static_aad_length[1196]       =   64'h0000000000000100;
assign   tb_i_aad[1196]                        =   tb_i_aad[1195];
assign   tb_i_rf_static_plaintext_length[1196] =   64'h0000000000000280;
assign   tb_i_plaintext[1196]                  =   tb_i_plaintext[1195];
assign   tb_o_valid[1196]                      =   1'b0;
assign   tb_o_sop[1196]                        =   1'b0;
assign   tb_o_ciphertext[1196]                 =   tb_o_ciphertext[1195];
assign   tb_o_tag_ready[1196]                  =   1'b0;
assign   tb_o_tag[1196]                        =   tb_o_tag[1195];

// CLK no. 1197/1240
// *************************************************
assign   tb_i_valid[1197]                      =   1'b0;
assign   tb_i_reset[1197]                      =   1'b0;
assign   tb_i_sop[1197]                        =   1'b0;
assign   tb_i_key_update[1197]                 =   1'b0;
assign   tb_i_key[1197]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1197]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1197]               =   1'b0;
assign   tb_i_rf_static_encrypt[1197]          =   1'b1;
assign   tb_i_clear_fault_flags[1197]          =   1'b0;
assign   tb_i_rf_static_aad_length[1197]       =   64'h0000000000000100;
assign   tb_i_aad[1197]                        =   tb_i_aad[1196];
assign   tb_i_rf_static_plaintext_length[1197] =   64'h0000000000000280;
assign   tb_i_plaintext[1197]                  =   tb_i_plaintext[1196];
assign   tb_o_valid[1197]                      =   1'b0;
assign   tb_o_sop[1197]                        =   1'b0;
assign   tb_o_ciphertext[1197]                 =   tb_o_ciphertext[1196];
assign   tb_o_tag_ready[1197]                  =   1'b0;
assign   tb_o_tag[1197]                        =   tb_o_tag[1196];

// CLK no. 1198/1240
// *************************************************
assign   tb_i_valid[1198]                      =   1'b0;
assign   tb_i_reset[1198]                      =   1'b0;
assign   tb_i_sop[1198]                        =   1'b0;
assign   tb_i_key_update[1198]                 =   1'b0;
assign   tb_i_key[1198]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1198]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1198]               =   1'b0;
assign   tb_i_rf_static_encrypt[1198]          =   1'b1;
assign   tb_i_clear_fault_flags[1198]          =   1'b0;
assign   tb_i_rf_static_aad_length[1198]       =   64'h0000000000000100;
assign   tb_i_aad[1198]                        =   tb_i_aad[1197];
assign   tb_i_rf_static_plaintext_length[1198] =   64'h0000000000000280;
assign   tb_i_plaintext[1198]                  =   tb_i_plaintext[1197];
assign   tb_o_valid[1198]                      =   1'b0;
assign   tb_o_sop[1198]                        =   1'b0;
assign   tb_o_ciphertext[1198]                 =   tb_o_ciphertext[1197];
assign   tb_o_tag_ready[1198]                  =   1'b0;
assign   tb_o_tag[1198]                        =   tb_o_tag[1197];

// CLK no. 1199/1240
// *************************************************
assign   tb_i_valid[1199]                      =   1'b0;
assign   tb_i_reset[1199]                      =   1'b0;
assign   tb_i_sop[1199]                        =   1'b0;
assign   tb_i_key_update[1199]                 =   1'b0;
assign   tb_i_key[1199]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1199]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1199]               =   1'b0;
assign   tb_i_rf_static_encrypt[1199]          =   1'b1;
assign   tb_i_clear_fault_flags[1199]          =   1'b0;
assign   tb_i_rf_static_aad_length[1199]       =   64'h0000000000000100;
assign   tb_i_aad[1199]                        =   tb_i_aad[1198];
assign   tb_i_rf_static_plaintext_length[1199] =   64'h0000000000000280;
assign   tb_i_plaintext[1199]                  =   tb_i_plaintext[1198];
assign   tb_o_valid[1199]                      =   1'b0;
assign   tb_o_sop[1199]                        =   1'b0;
assign   tb_o_ciphertext[1199]                 =   tb_o_ciphertext[1198];
assign   tb_o_tag_ready[1199]                  =   1'b0;
assign   tb_o_tag[1199]                        =   tb_o_tag[1198];

// CLK no. 1200/1240
// *************************************************
assign   tb_i_valid[1200]                      =   1'b0;
assign   tb_i_reset[1200]                      =   1'b0;
assign   tb_i_sop[1200]                        =   1'b0;
assign   tb_i_key_update[1200]                 =   1'b0;
assign   tb_i_key[1200]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1200]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1200]               =   1'b0;
assign   tb_i_rf_static_encrypt[1200]          =   1'b1;
assign   tb_i_clear_fault_flags[1200]          =   1'b0;
assign   tb_i_rf_static_aad_length[1200]       =   64'h0000000000000100;
assign   tb_i_aad[1200]                        =   tb_i_aad[1199];
assign   tb_i_rf_static_plaintext_length[1200] =   64'h0000000000000280;
assign   tb_i_plaintext[1200]                  =   tb_i_plaintext[1199];
assign   tb_o_valid[1200]                      =   1'b0;
assign   tb_o_sop[1200]                        =   1'b0;
assign   tb_o_ciphertext[1200]                 =   tb_o_ciphertext[1199];
assign   tb_o_tag_ready[1200]                  =   1'b0;
assign   tb_o_tag[1200]                        =   tb_o_tag[1199];

// CLK no. 1201/1240
// *************************************************
assign   tb_i_valid[1201]                      =   1'b0;
assign   tb_i_reset[1201]                      =   1'b0;
assign   tb_i_sop[1201]                        =   1'b0;
assign   tb_i_key_update[1201]                 =   1'b0;
assign   tb_i_key[1201]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1201]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1201]               =   1'b0;
assign   tb_i_rf_static_encrypt[1201]          =   1'b1;
assign   tb_i_clear_fault_flags[1201]          =   1'b0;
assign   tb_i_rf_static_aad_length[1201]       =   64'h0000000000000100;
assign   tb_i_aad[1201]                        =   tb_i_aad[1200];
assign   tb_i_rf_static_plaintext_length[1201] =   64'h0000000000000280;
assign   tb_i_plaintext[1201]                  =   tb_i_plaintext[1200];
assign   tb_o_valid[1201]                      =   1'b0;
assign   tb_o_sop[1201]                        =   1'b0;
assign   tb_o_ciphertext[1201]                 =   tb_o_ciphertext[1200];
assign   tb_o_tag_ready[1201]                  =   1'b0;
assign   tb_o_tag[1201]                        =   tb_o_tag[1200];

// CLK no. 1202/1240
// *************************************************
assign   tb_i_valid[1202]                      =   1'b0;
assign   tb_i_reset[1202]                      =   1'b0;
assign   tb_i_sop[1202]                        =   1'b0;
assign   tb_i_key_update[1202]                 =   1'b0;
assign   tb_i_key[1202]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1202]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1202]               =   1'b0;
assign   tb_i_rf_static_encrypt[1202]          =   1'b1;
assign   tb_i_clear_fault_flags[1202]          =   1'b0;
assign   tb_i_rf_static_aad_length[1202]       =   64'h0000000000000100;
assign   tb_i_aad[1202]                        =   tb_i_aad[1201];
assign   tb_i_rf_static_plaintext_length[1202] =   64'h0000000000000280;
assign   tb_i_plaintext[1202]                  =   tb_i_plaintext[1201];
assign   tb_o_valid[1202]                      =   1'b0;
assign   tb_o_sop[1202]                        =   1'b0;
assign   tb_o_ciphertext[1202]                 =   tb_o_ciphertext[1201];
assign   tb_o_tag_ready[1202]                  =   1'b0;
assign   tb_o_tag[1202]                        =   tb_o_tag[1201];

// CLK no. 1203/1240
// *************************************************
assign   tb_i_valid[1203]                      =   1'b0;
assign   tb_i_reset[1203]                      =   1'b0;
assign   tb_i_sop[1203]                        =   1'b0;
assign   tb_i_key_update[1203]                 =   1'b0;
assign   tb_i_key[1203]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1203]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1203]               =   1'b0;
assign   tb_i_rf_static_encrypt[1203]          =   1'b1;
assign   tb_i_clear_fault_flags[1203]          =   1'b0;
assign   tb_i_rf_static_aad_length[1203]       =   64'h0000000000000100;
assign   tb_i_aad[1203]                        =   tb_i_aad[1202];
assign   tb_i_rf_static_plaintext_length[1203] =   64'h0000000000000280;
assign   tb_i_plaintext[1203]                  =   tb_i_plaintext[1202];
assign   tb_o_valid[1203]                      =   1'b0;
assign   tb_o_sop[1203]                        =   1'b0;
assign   tb_o_ciphertext[1203]                 =   tb_o_ciphertext[1202];
assign   tb_o_tag_ready[1203]                  =   1'b0;
assign   tb_o_tag[1203]                        =   tb_o_tag[1202];

// CLK no. 1204/1240
// *************************************************
assign   tb_i_valid[1204]                      =   1'b0;
assign   tb_i_reset[1204]                      =   1'b0;
assign   tb_i_sop[1204]                        =   1'b0;
assign   tb_i_key_update[1204]                 =   1'b0;
assign   tb_i_key[1204]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1204]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1204]               =   1'b0;
assign   tb_i_rf_static_encrypt[1204]          =   1'b1;
assign   tb_i_clear_fault_flags[1204]          =   1'b0;
assign   tb_i_rf_static_aad_length[1204]       =   64'h0000000000000100;
assign   tb_i_aad[1204]                        =   tb_i_aad[1203];
assign   tb_i_rf_static_plaintext_length[1204] =   64'h0000000000000280;
assign   tb_i_plaintext[1204]                  =   tb_i_plaintext[1203];
assign   tb_o_valid[1204]                      =   1'b0;
assign   tb_o_sop[1204]                        =   1'b0;
assign   tb_o_ciphertext[1204]                 =   tb_o_ciphertext[1203];
assign   tb_o_tag_ready[1204]                  =   1'b0;
assign   tb_o_tag[1204]                        =   tb_o_tag[1203];

// CLK no. 1205/1240
// *************************************************
assign   tb_i_valid[1205]                      =   1'b0;
assign   tb_i_reset[1205]                      =   1'b0;
assign   tb_i_sop[1205]                        =   1'b0;
assign   tb_i_key_update[1205]                 =   1'b0;
assign   tb_i_key[1205]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1205]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1205]               =   1'b0;
assign   tb_i_rf_static_encrypt[1205]          =   1'b1;
assign   tb_i_clear_fault_flags[1205]          =   1'b0;
assign   tb_i_rf_static_aad_length[1205]       =   64'h0000000000000100;
assign   tb_i_aad[1205]                        =   tb_i_aad[1204];
assign   tb_i_rf_static_plaintext_length[1205] =   64'h0000000000000280;
assign   tb_i_plaintext[1205]                  =   tb_i_plaintext[1204];
assign   tb_o_valid[1205]                      =   1'b0;
assign   tb_o_sop[1205]                        =   1'b0;
assign   tb_o_ciphertext[1205]                 =   tb_o_ciphertext[1204];
assign   tb_o_tag_ready[1205]                  =   1'b0;
assign   tb_o_tag[1205]                        =   tb_o_tag[1204];

// CLK no. 1206/1240
// *************************************************
assign   tb_i_valid[1206]                      =   1'b0;
assign   tb_i_reset[1206]                      =   1'b0;
assign   tb_i_sop[1206]                        =   1'b0;
assign   tb_i_key_update[1206]                 =   1'b0;
assign   tb_i_key[1206]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1206]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1206]               =   1'b0;
assign   tb_i_rf_static_encrypt[1206]          =   1'b1;
assign   tb_i_clear_fault_flags[1206]          =   1'b0;
assign   tb_i_rf_static_aad_length[1206]       =   64'h0000000000000100;
assign   tb_i_aad[1206]                        =   tb_i_aad[1205];
assign   tb_i_rf_static_plaintext_length[1206] =   64'h0000000000000280;
assign   tb_i_plaintext[1206]                  =   tb_i_plaintext[1205];
assign   tb_o_valid[1206]                      =   1'b0;
assign   tb_o_sop[1206]                        =   1'b0;
assign   tb_o_ciphertext[1206]                 =   tb_o_ciphertext[1205];
assign   tb_o_tag_ready[1206]                  =   1'b0;
assign   tb_o_tag[1206]                        =   tb_o_tag[1205];

// CLK no. 1207/1240
// *************************************************
assign   tb_i_valid[1207]                      =   1'b0;
assign   tb_i_reset[1207]                      =   1'b0;
assign   tb_i_sop[1207]                        =   1'b0;
assign   tb_i_key_update[1207]                 =   1'b0;
assign   tb_i_key[1207]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1207]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1207]               =   1'b0;
assign   tb_i_rf_static_encrypt[1207]          =   1'b1;
assign   tb_i_clear_fault_flags[1207]          =   1'b0;
assign   tb_i_rf_static_aad_length[1207]       =   64'h0000000000000100;
assign   tb_i_aad[1207]                        =   tb_i_aad[1206];
assign   tb_i_rf_static_plaintext_length[1207] =   64'h0000000000000280;
assign   tb_i_plaintext[1207]                  =   tb_i_plaintext[1206];
assign   tb_o_valid[1207]                      =   1'b0;
assign   tb_o_sop[1207]                        =   1'b0;
assign   tb_o_ciphertext[1207]                 =   tb_o_ciphertext[1206];
assign   tb_o_tag_ready[1207]                  =   1'b0;
assign   tb_o_tag[1207]                        =   tb_o_tag[1206];

// CLK no. 1208/1240
// *************************************************
assign   tb_i_valid[1208]                      =   1'b0;
assign   tb_i_reset[1208]                      =   1'b0;
assign   tb_i_sop[1208]                        =   1'b0;
assign   tb_i_key_update[1208]                 =   1'b0;
assign   tb_i_key[1208]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1208]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1208]               =   1'b0;
assign   tb_i_rf_static_encrypt[1208]          =   1'b1;
assign   tb_i_clear_fault_flags[1208]          =   1'b0;
assign   tb_i_rf_static_aad_length[1208]       =   64'h0000000000000100;
assign   tb_i_aad[1208]                        =   tb_i_aad[1207];
assign   tb_i_rf_static_plaintext_length[1208] =   64'h0000000000000280;
assign   tb_i_plaintext[1208]                  =   tb_i_plaintext[1207];
assign   tb_o_valid[1208]                      =   1'b0;
assign   tb_o_sop[1208]                        =   1'b0;
assign   tb_o_ciphertext[1208]                 =   tb_o_ciphertext[1207];
assign   tb_o_tag_ready[1208]                  =   1'b0;
assign   tb_o_tag[1208]                        =   tb_o_tag[1207];

// CLK no. 1209/1240
// *************************************************
assign   tb_i_valid[1209]                      =   1'b0;
assign   tb_i_reset[1209]                      =   1'b0;
assign   tb_i_sop[1209]                        =   1'b0;
assign   tb_i_key_update[1209]                 =   1'b0;
assign   tb_i_key[1209]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1209]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1209]               =   1'b0;
assign   tb_i_rf_static_encrypt[1209]          =   1'b1;
assign   tb_i_clear_fault_flags[1209]          =   1'b0;
assign   tb_i_rf_static_aad_length[1209]       =   64'h0000000000000100;
assign   tb_i_aad[1209]                        =   tb_i_aad[1208];
assign   tb_i_rf_static_plaintext_length[1209] =   64'h0000000000000280;
assign   tb_i_plaintext[1209]                  =   tb_i_plaintext[1208];
assign   tb_o_valid[1209]                      =   1'b0;
assign   tb_o_sop[1209]                        =   1'b0;
assign   tb_o_ciphertext[1209]                 =   tb_o_ciphertext[1208];
assign   tb_o_tag_ready[1209]                  =   1'b0;
assign   tb_o_tag[1209]                        =   tb_o_tag[1208];

// CLK no. 1210/1240
// *************************************************
assign   tb_i_valid[1210]                      =   1'b0;
assign   tb_i_reset[1210]                      =   1'b0;
assign   tb_i_sop[1210]                        =   1'b0;
assign   tb_i_key_update[1210]                 =   1'b0;
assign   tb_i_key[1210]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1210]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1210]               =   1'b0;
assign   tb_i_rf_static_encrypt[1210]          =   1'b1;
assign   tb_i_clear_fault_flags[1210]          =   1'b0;
assign   tb_i_rf_static_aad_length[1210]       =   64'h0000000000000100;
assign   tb_i_aad[1210]                        =   tb_i_aad[1209];
assign   tb_i_rf_static_plaintext_length[1210] =   64'h0000000000000280;
assign   tb_i_plaintext[1210]                  =   tb_i_plaintext[1209];
assign   tb_o_valid[1210]                      =   1'b0;
assign   tb_o_sop[1210]                        =   1'b0;
assign   tb_o_ciphertext[1210]                 =   tb_o_ciphertext[1209];
assign   tb_o_tag_ready[1210]                  =   1'b0;
assign   tb_o_tag[1210]                        =   tb_o_tag[1209];

// CLK no. 1211/1240
// *************************************************
assign   tb_i_valid[1211]                      =   1'b0;
assign   tb_i_reset[1211]                      =   1'b0;
assign   tb_i_sop[1211]                        =   1'b0;
assign   tb_i_key_update[1211]                 =   1'b0;
assign   tb_i_key[1211]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1211]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1211]               =   1'b0;
assign   tb_i_rf_static_encrypt[1211]          =   1'b1;
assign   tb_i_clear_fault_flags[1211]          =   1'b0;
assign   tb_i_rf_static_aad_length[1211]       =   64'h0000000000000100;
assign   tb_i_aad[1211]                        =   tb_i_aad[1210];
assign   tb_i_rf_static_plaintext_length[1211] =   64'h0000000000000280;
assign   tb_i_plaintext[1211]                  =   tb_i_plaintext[1210];
assign   tb_o_valid[1211]                      =   1'b0;
assign   tb_o_sop[1211]                        =   1'b0;
assign   tb_o_ciphertext[1211]                 =   tb_o_ciphertext[1210];
assign   tb_o_tag_ready[1211]                  =   1'b0;
assign   tb_o_tag[1211]                        =   tb_o_tag[1210];

// CLK no. 1212/1240
// *************************************************
assign   tb_i_valid[1212]                      =   1'b0;
assign   tb_i_reset[1212]                      =   1'b0;
assign   tb_i_sop[1212]                        =   1'b0;
assign   tb_i_key_update[1212]                 =   1'b0;
assign   tb_i_key[1212]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1212]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1212]               =   1'b0;
assign   tb_i_rf_static_encrypt[1212]          =   1'b1;
assign   tb_i_clear_fault_flags[1212]          =   1'b0;
assign   tb_i_rf_static_aad_length[1212]       =   64'h0000000000000100;
assign   tb_i_aad[1212]                        =   tb_i_aad[1211];
assign   tb_i_rf_static_plaintext_length[1212] =   64'h0000000000000280;
assign   tb_i_plaintext[1212]                  =   tb_i_plaintext[1211];
assign   tb_o_valid[1212]                      =   1'b0;
assign   tb_o_sop[1212]                        =   1'b0;
assign   tb_o_ciphertext[1212]                 =   tb_o_ciphertext[1211];
assign   tb_o_tag_ready[1212]                  =   1'b0;
assign   tb_o_tag[1212]                        =   tb_o_tag[1211];

// CLK no. 1213/1240
// *************************************************
assign   tb_i_valid[1213]                      =   1'b0;
assign   tb_i_reset[1213]                      =   1'b0;
assign   tb_i_sop[1213]                        =   1'b0;
assign   tb_i_key_update[1213]                 =   1'b0;
assign   tb_i_key[1213]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1213]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1213]               =   1'b0;
assign   tb_i_rf_static_encrypt[1213]          =   1'b1;
assign   tb_i_clear_fault_flags[1213]          =   1'b0;
assign   tb_i_rf_static_aad_length[1213]       =   64'h0000000000000100;
assign   tb_i_aad[1213]                        =   tb_i_aad[1212];
assign   tb_i_rf_static_plaintext_length[1213] =   64'h0000000000000280;
assign   tb_i_plaintext[1213]                  =   tb_i_plaintext[1212];
assign   tb_o_valid[1213]                      =   1'b0;
assign   tb_o_sop[1213]                        =   1'b0;
assign   tb_o_ciphertext[1213]                 =   tb_o_ciphertext[1212];
assign   tb_o_tag_ready[1213]                  =   1'b0;
assign   tb_o_tag[1213]                        =   tb_o_tag[1212];

// CLK no. 1214/1240
// *************************************************
assign   tb_i_valid[1214]                      =   1'b0;
assign   tb_i_reset[1214]                      =   1'b0;
assign   tb_i_sop[1214]                        =   1'b0;
assign   tb_i_key_update[1214]                 =   1'b0;
assign   tb_i_key[1214]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1214]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1214]               =   1'b0;
assign   tb_i_rf_static_encrypt[1214]          =   1'b1;
assign   tb_i_clear_fault_flags[1214]          =   1'b0;
assign   tb_i_rf_static_aad_length[1214]       =   64'h0000000000000100;
assign   tb_i_aad[1214]                        =   tb_i_aad[1213];
assign   tb_i_rf_static_plaintext_length[1214] =   64'h0000000000000280;
assign   tb_i_plaintext[1214]                  =   tb_i_plaintext[1213];
assign   tb_o_valid[1214]                      =   1'b0;
assign   tb_o_sop[1214]                        =   1'b0;
assign   tb_o_ciphertext[1214]                 =   tb_o_ciphertext[1213];
assign   tb_o_tag_ready[1214]                  =   1'b0;
assign   tb_o_tag[1214]                        =   tb_o_tag[1213];

// CLK no. 1215/1240
// *************************************************
assign   tb_i_valid[1215]                      =   1'b0;
assign   tb_i_reset[1215]                      =   1'b0;
assign   tb_i_sop[1215]                        =   1'b0;
assign   tb_i_key_update[1215]                 =   1'b0;
assign   tb_i_key[1215]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1215]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1215]               =   1'b0;
assign   tb_i_rf_static_encrypt[1215]          =   1'b1;
assign   tb_i_clear_fault_flags[1215]          =   1'b0;
assign   tb_i_rf_static_aad_length[1215]       =   64'h0000000000000100;
assign   tb_i_aad[1215]                        =   tb_i_aad[1214];
assign   tb_i_rf_static_plaintext_length[1215] =   64'h0000000000000280;
assign   tb_i_plaintext[1215]                  =   tb_i_plaintext[1214];
assign   tb_o_valid[1215]                      =   1'b0;
assign   tb_o_sop[1215]                        =   1'b0;
assign   tb_o_ciphertext[1215]                 =   tb_o_ciphertext[1214];
assign   tb_o_tag_ready[1215]                  =   1'b0;
assign   tb_o_tag[1215]                        =   tb_o_tag[1214];

// CLK no. 1216/1240
// *************************************************
assign   tb_i_valid[1216]                      =   1'b0;
assign   tb_i_reset[1216]                      =   1'b0;
assign   tb_i_sop[1216]                        =   1'b0;
assign   tb_i_key_update[1216]                 =   1'b0;
assign   tb_i_key[1216]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1216]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1216]               =   1'b0;
assign   tb_i_rf_static_encrypt[1216]          =   1'b1;
assign   tb_i_clear_fault_flags[1216]          =   1'b0;
assign   tb_i_rf_static_aad_length[1216]       =   64'h0000000000000100;
assign   tb_i_aad[1216]                        =   tb_i_aad[1215];
assign   tb_i_rf_static_plaintext_length[1216] =   64'h0000000000000280;
assign   tb_i_plaintext[1216]                  =   tb_i_plaintext[1215];
assign   tb_o_valid[1216]                      =   1'b0;
assign   tb_o_sop[1216]                        =   1'b0;
assign   tb_o_ciphertext[1216]                 =   tb_o_ciphertext[1215];
assign   tb_o_tag_ready[1216]                  =   1'b0;
assign   tb_o_tag[1216]                        =   tb_o_tag[1215];

// CLK no. 1217/1240
// *************************************************
assign   tb_i_valid[1217]                      =   1'b0;
assign   tb_i_reset[1217]                      =   1'b0;
assign   tb_i_sop[1217]                        =   1'b0;
assign   tb_i_key_update[1217]                 =   1'b0;
assign   tb_i_key[1217]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1217]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1217]               =   1'b0;
assign   tb_i_rf_static_encrypt[1217]          =   1'b1;
assign   tb_i_clear_fault_flags[1217]          =   1'b0;
assign   tb_i_rf_static_aad_length[1217]       =   64'h0000000000000100;
assign   tb_i_aad[1217]                        =   tb_i_aad[1216];
assign   tb_i_rf_static_plaintext_length[1217] =   64'h0000000000000280;
assign   tb_i_plaintext[1217]                  =   tb_i_plaintext[1216];
assign   tb_o_valid[1217]                      =   1'b0;
assign   tb_o_sop[1217]                        =   1'b0;
assign   tb_o_ciphertext[1217]                 =   tb_o_ciphertext[1216];
assign   tb_o_tag_ready[1217]                  =   1'b0;
assign   tb_o_tag[1217]                        =   tb_o_tag[1216];

// CLK no. 1218/1240
// *************************************************
assign   tb_i_valid[1218]                      =   1'b0;
assign   tb_i_reset[1218]                      =   1'b0;
assign   tb_i_sop[1218]                        =   1'b0;
assign   tb_i_key_update[1218]                 =   1'b0;
assign   tb_i_key[1218]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1218]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1218]               =   1'b0;
assign   tb_i_rf_static_encrypt[1218]          =   1'b1;
assign   tb_i_clear_fault_flags[1218]          =   1'b0;
assign   tb_i_rf_static_aad_length[1218]       =   64'h0000000000000100;
assign   tb_i_aad[1218]                        =   tb_i_aad[1217];
assign   tb_i_rf_static_plaintext_length[1218] =   64'h0000000000000280;
assign   tb_i_plaintext[1218]                  =   tb_i_plaintext[1217];
assign   tb_o_valid[1218]                      =   1'b0;
assign   tb_o_sop[1218]                        =   1'b0;
assign   tb_o_ciphertext[1218]                 =   tb_o_ciphertext[1217];
assign   tb_o_tag_ready[1218]                  =   1'b0;
assign   tb_o_tag[1218]                        =   tb_o_tag[1217];

// CLK no. 1219/1240
// *************************************************
assign   tb_i_valid[1219]                      =   1'b0;
assign   tb_i_reset[1219]                      =   1'b0;
assign   tb_i_sop[1219]                        =   1'b0;
assign   tb_i_key_update[1219]                 =   1'b0;
assign   tb_i_key[1219]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1219]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1219]               =   1'b0;
assign   tb_i_rf_static_encrypt[1219]          =   1'b1;
assign   tb_i_clear_fault_flags[1219]          =   1'b0;
assign   tb_i_rf_static_aad_length[1219]       =   64'h0000000000000100;
assign   tb_i_aad[1219]                        =   tb_i_aad[1218];
assign   tb_i_rf_static_plaintext_length[1219] =   64'h0000000000000280;
assign   tb_i_plaintext[1219]                  =   tb_i_plaintext[1218];
assign   tb_o_valid[1219]                      =   1'b0;
assign   tb_o_sop[1219]                        =   1'b0;
assign   tb_o_ciphertext[1219]                 =   tb_o_ciphertext[1218];
assign   tb_o_tag_ready[1219]                  =   1'b0;
assign   tb_o_tag[1219]                        =   tb_o_tag[1218];

// CLK no. 1220/1240
// *************************************************
assign   tb_i_valid[1220]                      =   1'b0;
assign   tb_i_reset[1220]                      =   1'b0;
assign   tb_i_sop[1220]                        =   1'b0;
assign   tb_i_key_update[1220]                 =   1'b0;
assign   tb_i_key[1220]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1220]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1220]               =   1'b0;
assign   tb_i_rf_static_encrypt[1220]          =   1'b1;
assign   tb_i_clear_fault_flags[1220]          =   1'b0;
assign   tb_i_rf_static_aad_length[1220]       =   64'h0000000000000100;
assign   tb_i_aad[1220]                        =   tb_i_aad[1219];
assign   tb_i_rf_static_plaintext_length[1220] =   64'h0000000000000280;
assign   tb_i_plaintext[1220]                  =   tb_i_plaintext[1219];
assign   tb_o_valid[1220]                      =   1'b0;
assign   tb_o_sop[1220]                        =   1'b0;
assign   tb_o_ciphertext[1220]                 =   tb_o_ciphertext[1219];
assign   tb_o_tag_ready[1220]                  =   1'b0;
assign   tb_o_tag[1220]                        =   tb_o_tag[1219];

// CLK no. 1221/1240
// *************************************************
assign   tb_i_valid[1221]                      =   1'b0;
assign   tb_i_reset[1221]                      =   1'b0;
assign   tb_i_sop[1221]                        =   1'b0;
assign   tb_i_key_update[1221]                 =   1'b0;
assign   tb_i_key[1221]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1221]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1221]               =   1'b0;
assign   tb_i_rf_static_encrypt[1221]          =   1'b1;
assign   tb_i_clear_fault_flags[1221]          =   1'b0;
assign   tb_i_rf_static_aad_length[1221]       =   64'h0000000000000100;
assign   tb_i_aad[1221]                        =   tb_i_aad[1220];
assign   tb_i_rf_static_plaintext_length[1221] =   64'h0000000000000280;
assign   tb_i_plaintext[1221]                  =   tb_i_plaintext[1220];
assign   tb_o_valid[1221]                      =   1'b0;
assign   tb_o_sop[1221]                        =   1'b0;
assign   tb_o_ciphertext[1221]                 =   tb_o_ciphertext[1220];
assign   tb_o_tag_ready[1221]                  =   1'b0;
assign   tb_o_tag[1221]                        =   tb_o_tag[1220];

// CLK no. 1222/1240
// *************************************************
assign   tb_i_valid[1222]                      =   1'b0;
assign   tb_i_reset[1222]                      =   1'b0;
assign   tb_i_sop[1222]                        =   1'b0;
assign   tb_i_key_update[1222]                 =   1'b0;
assign   tb_i_key[1222]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1222]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1222]               =   1'b0;
assign   tb_i_rf_static_encrypt[1222]          =   1'b1;
assign   tb_i_clear_fault_flags[1222]          =   1'b0;
assign   tb_i_rf_static_aad_length[1222]       =   64'h0000000000000100;
assign   tb_i_aad[1222]                        =   tb_i_aad[1221];
assign   tb_i_rf_static_plaintext_length[1222] =   64'h0000000000000280;
assign   tb_i_plaintext[1222]                  =   tb_i_plaintext[1221];
assign   tb_o_valid[1222]                      =   1'b0;
assign   tb_o_sop[1222]                        =   1'b0;
assign   tb_o_ciphertext[1222]                 =   tb_o_ciphertext[1221];
assign   tb_o_tag_ready[1222]                  =   1'b0;
assign   tb_o_tag[1222]                        =   tb_o_tag[1221];

// CLK no. 1223/1240
// *************************************************
assign   tb_i_valid[1223]                      =   1'b0;
assign   tb_i_reset[1223]                      =   1'b0;
assign   tb_i_sop[1223]                        =   1'b0;
assign   tb_i_key_update[1223]                 =   1'b0;
assign   tb_i_key[1223]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1223]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1223]               =   1'b0;
assign   tb_i_rf_static_encrypt[1223]          =   1'b1;
assign   tb_i_clear_fault_flags[1223]          =   1'b0;
assign   tb_i_rf_static_aad_length[1223]       =   64'h0000000000000100;
assign   tb_i_aad[1223]                        =   tb_i_aad[1222];
assign   tb_i_rf_static_plaintext_length[1223] =   64'h0000000000000280;
assign   tb_i_plaintext[1223]                  =   tb_i_plaintext[1222];
assign   tb_o_valid[1223]                      =   1'b0;
assign   tb_o_sop[1223]                        =   1'b0;
assign   tb_o_ciphertext[1223]                 =   tb_o_ciphertext[1222];
assign   tb_o_tag_ready[1223]                  =   1'b0;
assign   tb_o_tag[1223]                        =   tb_o_tag[1222];

// CLK no. 1224/1240
// *************************************************
assign   tb_i_valid[1224]                      =   1'b0;
assign   tb_i_reset[1224]                      =   1'b0;
assign   tb_i_sop[1224]                        =   1'b0;
assign   tb_i_key_update[1224]                 =   1'b0;
assign   tb_i_key[1224]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1224]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1224]               =   1'b0;
assign   tb_i_rf_static_encrypt[1224]          =   1'b1;
assign   tb_i_clear_fault_flags[1224]          =   1'b0;
assign   tb_i_rf_static_aad_length[1224]       =   64'h0000000000000100;
assign   tb_i_aad[1224]                        =   tb_i_aad[1223];
assign   tb_i_rf_static_plaintext_length[1224] =   64'h0000000000000280;
assign   tb_i_plaintext[1224]                  =   tb_i_plaintext[1223];
assign   tb_o_valid[1224]                      =   1'b0;
assign   tb_o_sop[1224]                        =   1'b0;
assign   tb_o_ciphertext[1224]                 =   tb_o_ciphertext[1223];
assign   tb_o_tag_ready[1224]                  =   1'b0;
assign   tb_o_tag[1224]                        =   tb_o_tag[1223];

// CLK no. 1225/1240
// *************************************************
assign   tb_i_valid[1225]                      =   1'b0;
assign   tb_i_reset[1225]                      =   1'b0;
assign   tb_i_sop[1225]                        =   1'b0;
assign   tb_i_key_update[1225]                 =   1'b0;
assign   tb_i_key[1225]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1225]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1225]               =   1'b0;
assign   tb_i_rf_static_encrypt[1225]          =   1'b1;
assign   tb_i_clear_fault_flags[1225]          =   1'b0;
assign   tb_i_rf_static_aad_length[1225]       =   64'h0000000000000100;
assign   tb_i_aad[1225]                        =   tb_i_aad[1224];
assign   tb_i_rf_static_plaintext_length[1225] =   64'h0000000000000280;
assign   tb_i_plaintext[1225]                  =   tb_i_plaintext[1224];
assign   tb_o_valid[1225]                      =   1'b0;
assign   tb_o_sop[1225]                        =   1'b0;
assign   tb_o_ciphertext[1225]                 =   tb_o_ciphertext[1224];
assign   tb_o_tag_ready[1225]                  =   1'b0;
assign   tb_o_tag[1225]                        =   tb_o_tag[1224];

// CLK no. 1226/1240
// *************************************************
assign   tb_i_valid[1226]                      =   1'b0;
assign   tb_i_reset[1226]                      =   1'b0;
assign   tb_i_sop[1226]                        =   1'b0;
assign   tb_i_key_update[1226]                 =   1'b0;
assign   tb_i_key[1226]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1226]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1226]               =   1'b0;
assign   tb_i_rf_static_encrypt[1226]          =   1'b1;
assign   tb_i_clear_fault_flags[1226]          =   1'b0;
assign   tb_i_rf_static_aad_length[1226]       =   64'h0000000000000100;
assign   tb_i_aad[1226]                        =   tb_i_aad[1225];
assign   tb_i_rf_static_plaintext_length[1226] =   64'h0000000000000280;
assign   tb_i_plaintext[1226]                  =   tb_i_plaintext[1225];
assign   tb_o_valid[1226]                      =   1'b0;
assign   tb_o_sop[1226]                        =   1'b0;
assign   tb_o_ciphertext[1226]                 =   tb_o_ciphertext[1225];
assign   tb_o_tag_ready[1226]                  =   1'b0;
assign   tb_o_tag[1226]                        =   tb_o_tag[1225];

// CLK no. 1227/1240
// *************************************************
assign   tb_i_valid[1227]                      =   1'b0;
assign   tb_i_reset[1227]                      =   1'b0;
assign   tb_i_sop[1227]                        =   1'b0;
assign   tb_i_key_update[1227]                 =   1'b0;
assign   tb_i_key[1227]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1227]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1227]               =   1'b0;
assign   tb_i_rf_static_encrypt[1227]          =   1'b1;
assign   tb_i_clear_fault_flags[1227]          =   1'b0;
assign   tb_i_rf_static_aad_length[1227]       =   64'h0000000000000100;
assign   tb_i_aad[1227]                        =   tb_i_aad[1226];
assign   tb_i_rf_static_plaintext_length[1227] =   64'h0000000000000280;
assign   tb_i_plaintext[1227]                  =   tb_i_plaintext[1226];
assign   tb_o_valid[1227]                      =   1'b1;
assign   tb_o_sop[1227]                        =   1'b1;
assign   tb_o_ciphertext[1227]                 =   256'hae37ed45d6c795509dbbb4bdec9d6b730aeb19372444786c589db791d5c87242;
assign   tb_o_tag_ready[1227]                  =   1'b0;
assign   tb_o_tag[1227]                        =   tb_o_tag[1226];

// CLK no. 1228/1240
// *************************************************
assign   tb_i_valid[1228]                      =   1'b0;
assign   tb_i_reset[1228]                      =   1'b0;
assign   tb_i_sop[1228]                        =   1'b0;
assign   tb_i_key_update[1228]                 =   1'b0;
assign   tb_i_key[1228]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1228]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1228]               =   1'b0;
assign   tb_i_rf_static_encrypt[1228]          =   1'b1;
assign   tb_i_clear_fault_flags[1228]          =   1'b0;
assign   tb_i_rf_static_aad_length[1228]       =   64'h0000000000000100;
assign   tb_i_aad[1228]                        =   tb_i_aad[1227];
assign   tb_i_rf_static_plaintext_length[1228] =   64'h0000000000000280;
assign   tb_i_plaintext[1228]                  =   tb_i_plaintext[1227];
assign   tb_o_valid[1228]                      =   1'b1;
assign   tb_o_sop[1228]                        =   1'b0;
assign   tb_o_ciphertext[1228]                 =   256'h9b4a55e0081e65324b941027d9fc9520edb58e64a928b84694997a277f08ae9d;
assign   tb_o_tag_ready[1228]                  =   1'b0;
assign   tb_o_tag[1228]                        =   tb_o_tag[1227];

// CLK no. 1229/1240
// *************************************************
assign   tb_i_valid[1229]                      =   1'b0;
assign   tb_i_reset[1229]                      =   1'b0;
assign   tb_i_sop[1229]                        =   1'b0;
assign   tb_i_key_update[1229]                 =   1'b0;
assign   tb_i_key[1229]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1229]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1229]               =   1'b0;
assign   tb_i_rf_static_encrypt[1229]          =   1'b1;
assign   tb_i_clear_fault_flags[1229]          =   1'b0;
assign   tb_i_rf_static_aad_length[1229]       =   64'h0000000000000100;
assign   tb_i_aad[1229]                        =   tb_i_aad[1228];
assign   tb_i_rf_static_plaintext_length[1229] =   64'h0000000000000280;
assign   tb_i_plaintext[1229]                  =   tb_i_plaintext[1228];
assign   tb_o_valid[1229]                      =   1'b1;
assign   tb_o_sop[1229]                        =   1'b0;
assign   tb_o_ciphertext[1229]                 =   256'h332d0a43e9980d5b2090d02a549a2ab9;
assign   tb_o_tag_ready[1229]                  =   1'b0;
assign   tb_o_tag[1229]                        =   tb_o_tag[1228];

// CLK no. 1230/1240
// *************************************************
assign   tb_i_valid[1230]                      =   1'b0;
assign   tb_i_reset[1230]                      =   1'b0;
assign   tb_i_sop[1230]                        =   1'b0;
assign   tb_i_key_update[1230]                 =   1'b0;
assign   tb_i_key[1230]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1230]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1230]               =   1'b0;
assign   tb_i_rf_static_encrypt[1230]          =   1'b1;
assign   tb_i_clear_fault_flags[1230]          =   1'b0;
assign   tb_i_rf_static_aad_length[1230]       =   64'h0000000000000100;
assign   tb_i_aad[1230]                        =   tb_i_aad[1229];
assign   tb_i_rf_static_plaintext_length[1230] =   64'h0000000000000280;
assign   tb_i_plaintext[1230]                  =   tb_i_plaintext[1229];
assign   tb_o_valid[1230]                      =   1'b0;
assign   tb_o_sop[1230]                        =   1'b0;
assign   tb_o_ciphertext[1230]                 =   tb_o_ciphertext[1229];
assign   tb_o_tag_ready[1230]                  =   1'b0;
assign   tb_o_tag[1230]                        =   tb_o_tag[1229];

// CLK no. 1231/1240
// *************************************************
assign   tb_i_valid[1231]                      =   1'b0;
assign   tb_i_reset[1231]                      =   1'b0;
assign   tb_i_sop[1231]                        =   1'b0;
assign   tb_i_key_update[1231]                 =   1'b0;
assign   tb_i_key[1231]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1231]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1231]               =   1'b0;
assign   tb_i_rf_static_encrypt[1231]          =   1'b1;
assign   tb_i_clear_fault_flags[1231]          =   1'b0;
assign   tb_i_rf_static_aad_length[1231]       =   64'h0000000000000100;
assign   tb_i_aad[1231]                        =   tb_i_aad[1230];
assign   tb_i_rf_static_plaintext_length[1231] =   64'h0000000000000280;
assign   tb_i_plaintext[1231]                  =   tb_i_plaintext[1230];
assign   tb_o_valid[1231]                      =   1'b0;
assign   tb_o_sop[1231]                        =   1'b0;
assign   tb_o_ciphertext[1231]                 =   tb_o_ciphertext[1230];
assign   tb_o_tag_ready[1231]                  =   1'b0;
assign   tb_o_tag[1231]                        =   tb_o_tag[1230];

// CLK no. 1232/1240
// *************************************************
assign   tb_i_valid[1232]                      =   1'b0;
assign   tb_i_reset[1232]                      =   1'b0;
assign   tb_i_sop[1232]                        =   1'b0;
assign   tb_i_key_update[1232]                 =   1'b0;
assign   tb_i_key[1232]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1232]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1232]               =   1'b0;
assign   tb_i_rf_static_encrypt[1232]          =   1'b1;
assign   tb_i_clear_fault_flags[1232]          =   1'b0;
assign   tb_i_rf_static_aad_length[1232]       =   64'h0000000000000100;
assign   tb_i_aad[1232]                        =   tb_i_aad[1231];
assign   tb_i_rf_static_plaintext_length[1232] =   64'h0000000000000280;
assign   tb_i_plaintext[1232]                  =   tb_i_plaintext[1231];
assign   tb_o_valid[1232]                      =   1'b0;
assign   tb_o_sop[1232]                        =   1'b0;
assign   tb_o_ciphertext[1232]                 =   tb_o_ciphertext[1231];
assign   tb_o_tag_ready[1232]                  =   1'b0;
assign   tb_o_tag[1232]                        =   tb_o_tag[1231];

// CLK no. 1233/1240
// *************************************************
assign   tb_i_valid[1233]                      =   1'b0;
assign   tb_i_reset[1233]                      =   1'b0;
assign   tb_i_sop[1233]                        =   1'b0;
assign   tb_i_key_update[1233]                 =   1'b0;
assign   tb_i_key[1233]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1233]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1233]               =   1'b0;
assign   tb_i_rf_static_encrypt[1233]          =   1'b1;
assign   tb_i_clear_fault_flags[1233]          =   1'b0;
assign   tb_i_rf_static_aad_length[1233]       =   64'h0000000000000100;
assign   tb_i_aad[1233]                        =   tb_i_aad[1232];
assign   tb_i_rf_static_plaintext_length[1233] =   64'h0000000000000280;
assign   tb_i_plaintext[1233]                  =   tb_i_plaintext[1232];
assign   tb_o_valid[1233]                      =   1'b0;
assign   tb_o_sop[1233]                        =   1'b0;
assign   tb_o_ciphertext[1233]                 =   tb_o_ciphertext[1232];
assign   tb_o_tag_ready[1233]                  =   1'b0;
assign   tb_o_tag[1233]                        =   tb_o_tag[1232];

// CLK no. 1234/1240
// *************************************************
assign   tb_i_valid[1234]                      =   1'b0;
assign   tb_i_reset[1234]                      =   1'b0;
assign   tb_i_sop[1234]                        =   1'b0;
assign   tb_i_key_update[1234]                 =   1'b0;
assign   tb_i_key[1234]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1234]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1234]               =   1'b0;
assign   tb_i_rf_static_encrypt[1234]          =   1'b1;
assign   tb_i_clear_fault_flags[1234]          =   1'b0;
assign   tb_i_rf_static_aad_length[1234]       =   64'h0000000000000100;
assign   tb_i_aad[1234]                        =   tb_i_aad[1233];
assign   tb_i_rf_static_plaintext_length[1234] =   64'h0000000000000280;
assign   tb_i_plaintext[1234]                  =   tb_i_plaintext[1233];
assign   tb_o_valid[1234]                      =   1'b0;
assign   tb_o_sop[1234]                        =   1'b0;
assign   tb_o_ciphertext[1234]                 =   tb_o_ciphertext[1233];
assign   tb_o_tag_ready[1234]                  =   1'b0;
assign   tb_o_tag[1234]                        =   tb_o_tag[1233];

// CLK no. 1235/1240
// *************************************************
assign   tb_i_valid[1235]                      =   1'b0;
assign   tb_i_reset[1235]                      =   1'b0;
assign   tb_i_sop[1235]                        =   1'b0;
assign   tb_i_key_update[1235]                 =   1'b0;
assign   tb_i_key[1235]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1235]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1235]               =   1'b0;
assign   tb_i_rf_static_encrypt[1235]          =   1'b1;
assign   tb_i_clear_fault_flags[1235]          =   1'b0;
assign   tb_i_rf_static_aad_length[1235]       =   64'h0000000000000100;
assign   tb_i_aad[1235]                        =   tb_i_aad[1234];
assign   tb_i_rf_static_plaintext_length[1235] =   64'h0000000000000280;
assign   tb_i_plaintext[1235]                  =   tb_i_plaintext[1234];
assign   tb_o_valid[1235]                      =   1'b0;
assign   tb_o_sop[1235]                        =   1'b0;
assign   tb_o_ciphertext[1235]                 =   tb_o_ciphertext[1234];
assign   tb_o_tag_ready[1235]                  =   1'b0;
assign   tb_o_tag[1235]                        =   tb_o_tag[1234];

// CLK no. 1236/1240
// *************************************************
assign   tb_i_valid[1236]                      =   1'b0;
assign   tb_i_reset[1236]                      =   1'b0;
assign   tb_i_sop[1236]                        =   1'b0;
assign   tb_i_key_update[1236]                 =   1'b0;
assign   tb_i_key[1236]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1236]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1236]               =   1'b0;
assign   tb_i_rf_static_encrypt[1236]          =   1'b1;
assign   tb_i_clear_fault_flags[1236]          =   1'b0;
assign   tb_i_rf_static_aad_length[1236]       =   64'h0000000000000100;
assign   tb_i_aad[1236]                        =   tb_i_aad[1235];
assign   tb_i_rf_static_plaintext_length[1236] =   64'h0000000000000280;
assign   tb_i_plaintext[1236]                  =   tb_i_plaintext[1235];
assign   tb_o_valid[1236]                      =   1'b0;
assign   tb_o_sop[1236]                        =   1'b0;
assign   tb_o_ciphertext[1236]                 =   tb_o_ciphertext[1235];
assign   tb_o_tag_ready[1236]                  =   1'b0;
assign   tb_o_tag[1236]                        =   tb_o_tag[1235];

// CLK no. 1237/1240
// *************************************************
assign   tb_i_valid[1237]                      =   1'b0;
assign   tb_i_reset[1237]                      =   1'b0;
assign   tb_i_sop[1237]                        =   1'b0;
assign   tb_i_key_update[1237]                 =   1'b0;
assign   tb_i_key[1237]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1237]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1237]               =   1'b0;
assign   tb_i_rf_static_encrypt[1237]          =   1'b1;
assign   tb_i_clear_fault_flags[1237]          =   1'b0;
assign   tb_i_rf_static_aad_length[1237]       =   64'h0000000000000100;
assign   tb_i_aad[1237]                        =   tb_i_aad[1236];
assign   tb_i_rf_static_plaintext_length[1237] =   64'h0000000000000280;
assign   tb_i_plaintext[1237]                  =   tb_i_plaintext[1236];
assign   tb_o_valid[1237]                      =   1'b0;
assign   tb_o_sop[1237]                        =   1'b0;
assign   tb_o_ciphertext[1237]                 =   tb_o_ciphertext[1236];
assign   tb_o_tag_ready[1237]                  =   1'b1;
assign   tb_o_tag[1237]                        =   128'h5d34a0f4221bc8300c3bbe8ace3cd548;

// CLK no. 1238/1240
// *************************************************
assign   tb_i_valid[1238]                      =   1'b0;
assign   tb_i_reset[1238]                      =   1'b0;
assign   tb_i_sop[1238]                        =   1'b0;
assign   tb_i_key_update[1238]                 =   1'b0;
assign   tb_i_key[1238]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1238]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1238]               =   1'b0;
assign   tb_i_rf_static_encrypt[1238]          =   1'b1;
assign   tb_i_clear_fault_flags[1238]          =   1'b0;
assign   tb_i_rf_static_aad_length[1238]       =   64'h0000000000000100;
assign   tb_i_aad[1238]                        =   tb_i_aad[1237];
assign   tb_i_rf_static_plaintext_length[1238] =   64'h0000000000000280;
assign   tb_i_plaintext[1238]                  =   tb_i_plaintext[1237];
assign   tb_o_valid[1238]                      =   1'b0;
assign   tb_o_sop[1238]                        =   1'b0;
assign   tb_o_ciphertext[1238]                 =   tb_o_ciphertext[1237];
assign   tb_o_tag_ready[1238]                  =   1'b0;
assign   tb_o_tag[1238]                        =   tb_o_tag[1237];

// CLK no. 1239/1240
// *************************************************
assign   tb_i_valid[1239]                      =   1'b0;
assign   tb_i_reset[1239]                      =   1'b0;
assign   tb_i_sop[1239]                        =   1'b0;
assign   tb_i_key_update[1239]                 =   1'b0;
assign   tb_i_key[1239]                        =   256'hfeffe9928665731c6d6a8f9467308308feffe9928665731c6d6a8f9467308308;
assign   tb_i_iv[1239]                         =   96'hcafebabefacedbaddecaf888;
assign   tb_i_rf_mode_gmac[1239]               =   1'b0;
assign   tb_i_rf_static_encrypt[1239]          =   1'b1;
assign   tb_i_clear_fault_flags[1239]          =   1'b0;
assign   tb_i_rf_static_aad_length[1239]       =   64'h0000000000000100;
assign   tb_i_aad[1239]                        =   tb_i_aad[1238];
assign   tb_i_rf_static_plaintext_length[1239] =   64'h0000000000000280;
assign   tb_i_plaintext[1239]                  =   tb_i_plaintext[1238];
assign   tb_o_valid[1239]                      =   1'b0;
assign   tb_o_sop[1239]                        =   1'b0;
assign   tb_o_ciphertext[1239]                 =   tb_o_ciphertext[1238];
assign   tb_o_tag_ready[1239]                  =   1'b0;
assign   tb_o_tag[1239]                        =   tb_o_tag[1238];

endmodule